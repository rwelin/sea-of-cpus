
library ieee;
use ieee.std_logic_1164.all;
use work.core_config.all;
use work.all;

entity Grid8x8 is
    port (
        clk: in std_logic;
        clk_en: in std_logic;
        reset: in std_logic;
        addr: in ram_addr;
        data: in word;
        we: in std_logic;
        fifo_inputs: in core_fifo_inputs_t;
        fifo_full: out std_logic_vector(0 to NUM_CORE_FIFOS-1);
        outputs: out core_fifo_inputs_t;
        outputs_full: in std_logic_vector(0 to NUM_CORE_FIFOS-1)
    );
end Grid8x8;

architecture behav of Grid8x8 is

    
        signal fifo_inputs_140095589890200: core_fifo_inputs_t;
        signal fifo_full_140095589890200: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589890200: core_fifo_inputs_t;
        signal outputs_full_140095589890200: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589890424: core_fifo_inputs_t;
        signal fifo_full_140095589890424: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589890424: core_fifo_inputs_t;
        signal outputs_full_140095589890424: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589890368: core_fifo_inputs_t;
        signal fifo_full_140095589890368: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589890368: core_fifo_inputs_t;
        signal outputs_full_140095589890368: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589890480: core_fifo_inputs_t;
        signal fifo_full_140095589890480: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589890480: core_fifo_inputs_t;
        signal outputs_full_140095589890480: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589890536: core_fifo_inputs_t;
        signal fifo_full_140095589890536: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589890536: core_fifo_inputs_t;
        signal outputs_full_140095589890536: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589890592: core_fifo_inputs_t;
        signal fifo_full_140095589890592: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589890592: core_fifo_inputs_t;
        signal outputs_full_140095589890592: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589890648: core_fifo_inputs_t;
        signal fifo_full_140095589890648: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589890648: core_fifo_inputs_t;
        signal outputs_full_140095589890648: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589890704: core_fifo_inputs_t;
        signal fifo_full_140095589890704: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589890704: core_fifo_inputs_t;
        signal outputs_full_140095589890704: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589890760: core_fifo_inputs_t;
        signal fifo_full_140095589890760: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589890760: core_fifo_inputs_t;
        signal outputs_full_140095589890760: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589890312: core_fifo_inputs_t;
        signal fifo_full_140095589890312: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589890312: core_fifo_inputs_t;
        signal outputs_full_140095589890312: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589890816: core_fifo_inputs_t;
        signal fifo_full_140095589890816: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589890816: core_fifo_inputs_t;
        signal outputs_full_140095589890816: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589890872: core_fifo_inputs_t;
        signal fifo_full_140095589890872: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589890872: core_fifo_inputs_t;
        signal outputs_full_140095589890872: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589890928: core_fifo_inputs_t;
        signal fifo_full_140095589890928: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589890928: core_fifo_inputs_t;
        signal outputs_full_140095589890928: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589890984: core_fifo_inputs_t;
        signal fifo_full_140095589890984: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589890984: core_fifo_inputs_t;
        signal outputs_full_140095589890984: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589891040: core_fifo_inputs_t;
        signal fifo_full_140095589891040: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589891040: core_fifo_inputs_t;
        signal outputs_full_140095589891040: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589891096: core_fifo_inputs_t;
        signal fifo_full_140095589891096: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589891096: core_fifo_inputs_t;
        signal outputs_full_140095589891096: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589891152: core_fifo_inputs_t;
        signal fifo_full_140095589891152: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589891152: core_fifo_inputs_t;
        signal outputs_full_140095589891152: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589891208: core_fifo_inputs_t;
        signal fifo_full_140095589891208: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589891208: core_fifo_inputs_t;
        signal outputs_full_140095589891208: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589891264: core_fifo_inputs_t;
        signal fifo_full_140095589891264: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589891264: core_fifo_inputs_t;
        signal outputs_full_140095589891264: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589891320: core_fifo_inputs_t;
        signal fifo_full_140095589891320: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589891320: core_fifo_inputs_t;
        signal outputs_full_140095589891320: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589891376: core_fifo_inputs_t;
        signal fifo_full_140095589891376: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589891376: core_fifo_inputs_t;
        signal outputs_full_140095589891376: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589891432: core_fifo_inputs_t;
        signal fifo_full_140095589891432: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589891432: core_fifo_inputs_t;
        signal outputs_full_140095589891432: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589891488: core_fifo_inputs_t;
        signal fifo_full_140095589891488: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589891488: core_fifo_inputs_t;
        signal outputs_full_140095589891488: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589891544: core_fifo_inputs_t;
        signal fifo_full_140095589891544: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589891544: core_fifo_inputs_t;
        signal outputs_full_140095589891544: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589891600: core_fifo_inputs_t;
        signal fifo_full_140095589891600: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589891600: core_fifo_inputs_t;
        signal outputs_full_140095589891600: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589891656: core_fifo_inputs_t;
        signal fifo_full_140095589891656: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589891656: core_fifo_inputs_t;
        signal outputs_full_140095589891656: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589891712: core_fifo_inputs_t;
        signal fifo_full_140095589891712: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589891712: core_fifo_inputs_t;
        signal outputs_full_140095589891712: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589891768: core_fifo_inputs_t;
        signal fifo_full_140095589891768: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589891768: core_fifo_inputs_t;
        signal outputs_full_140095589891768: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589891824: core_fifo_inputs_t;
        signal fifo_full_140095589891824: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589891824: core_fifo_inputs_t;
        signal outputs_full_140095589891824: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589891880: core_fifo_inputs_t;
        signal fifo_full_140095589891880: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589891880: core_fifo_inputs_t;
        signal outputs_full_140095589891880: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589891936: core_fifo_inputs_t;
        signal fifo_full_140095589891936: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589891936: core_fifo_inputs_t;
        signal outputs_full_140095589891936: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589891992: core_fifo_inputs_t;
        signal fifo_full_140095589891992: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589891992: core_fifo_inputs_t;
        signal outputs_full_140095589891992: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589892048: core_fifo_inputs_t;
        signal fifo_full_140095589892048: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589892048: core_fifo_inputs_t;
        signal outputs_full_140095589892048: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589933128: core_fifo_inputs_t;
        signal fifo_full_140095589933128: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589933128: core_fifo_inputs_t;
        signal outputs_full_140095589933128: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589933184: core_fifo_inputs_t;
        signal fifo_full_140095589933184: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589933184: core_fifo_inputs_t;
        signal outputs_full_140095589933184: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589933240: core_fifo_inputs_t;
        signal fifo_full_140095589933240: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589933240: core_fifo_inputs_t;
        signal outputs_full_140095589933240: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589933296: core_fifo_inputs_t;
        signal fifo_full_140095589933296: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589933296: core_fifo_inputs_t;
        signal outputs_full_140095589933296: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589933352: core_fifo_inputs_t;
        signal fifo_full_140095589933352: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589933352: core_fifo_inputs_t;
        signal outputs_full_140095589933352: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589933408: core_fifo_inputs_t;
        signal fifo_full_140095589933408: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589933408: core_fifo_inputs_t;
        signal outputs_full_140095589933408: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589933464: core_fifo_inputs_t;
        signal fifo_full_140095589933464: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589933464: core_fifo_inputs_t;
        signal outputs_full_140095589933464: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589933520: core_fifo_inputs_t;
        signal fifo_full_140095589933520: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589933520: core_fifo_inputs_t;
        signal outputs_full_140095589933520: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589933576: core_fifo_inputs_t;
        signal fifo_full_140095589933576: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589933576: core_fifo_inputs_t;
        signal outputs_full_140095589933576: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589933632: core_fifo_inputs_t;
        signal fifo_full_140095589933632: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589933632: core_fifo_inputs_t;
        signal outputs_full_140095589933632: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589933688: core_fifo_inputs_t;
        signal fifo_full_140095589933688: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589933688: core_fifo_inputs_t;
        signal outputs_full_140095589933688: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589933744: core_fifo_inputs_t;
        signal fifo_full_140095589933744: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589933744: core_fifo_inputs_t;
        signal outputs_full_140095589933744: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589933800: core_fifo_inputs_t;
        signal fifo_full_140095589933800: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589933800: core_fifo_inputs_t;
        signal outputs_full_140095589933800: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589933856: core_fifo_inputs_t;
        signal fifo_full_140095589933856: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589933856: core_fifo_inputs_t;
        signal outputs_full_140095589933856: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589933912: core_fifo_inputs_t;
        signal fifo_full_140095589933912: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589933912: core_fifo_inputs_t;
        signal outputs_full_140095589933912: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589933968: core_fifo_inputs_t;
        signal fifo_full_140095589933968: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589933968: core_fifo_inputs_t;
        signal outputs_full_140095589933968: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589934024: core_fifo_inputs_t;
        signal fifo_full_140095589934024: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589934024: core_fifo_inputs_t;
        signal outputs_full_140095589934024: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589934080: core_fifo_inputs_t;
        signal fifo_full_140095589934080: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589934080: core_fifo_inputs_t;
        signal outputs_full_140095589934080: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589934136: core_fifo_inputs_t;
        signal fifo_full_140095589934136: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589934136: core_fifo_inputs_t;
        signal outputs_full_140095589934136: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589934192: core_fifo_inputs_t;
        signal fifo_full_140095589934192: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589934192: core_fifo_inputs_t;
        signal outputs_full_140095589934192: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589934248: core_fifo_inputs_t;
        signal fifo_full_140095589934248: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589934248: core_fifo_inputs_t;
        signal outputs_full_140095589934248: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589934304: core_fifo_inputs_t;
        signal fifo_full_140095589934304: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589934304: core_fifo_inputs_t;
        signal outputs_full_140095589934304: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589934360: core_fifo_inputs_t;
        signal fifo_full_140095589934360: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589934360: core_fifo_inputs_t;
        signal outputs_full_140095589934360: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589934416: core_fifo_inputs_t;
        signal fifo_full_140095589934416: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589934416: core_fifo_inputs_t;
        signal outputs_full_140095589934416: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589934472: core_fifo_inputs_t;
        signal fifo_full_140095589934472: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589934472: core_fifo_inputs_t;
        signal outputs_full_140095589934472: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589934528: core_fifo_inputs_t;
        signal fifo_full_140095589934528: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589934528: core_fifo_inputs_t;
        signal outputs_full_140095589934528: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589934584: core_fifo_inputs_t;
        signal fifo_full_140095589934584: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589934584: core_fifo_inputs_t;
        signal outputs_full_140095589934584: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589934640: core_fifo_inputs_t;
        signal fifo_full_140095589934640: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589934640: core_fifo_inputs_t;
        signal outputs_full_140095589934640: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589934696: core_fifo_inputs_t;
        signal fifo_full_140095589934696: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589934696: core_fifo_inputs_t;
        signal outputs_full_140095589934696: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589934752: core_fifo_inputs_t;
        signal fifo_full_140095589934752: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589934752: core_fifo_inputs_t;
        signal outputs_full_140095589934752: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140095589934808: core_fifo_inputs_t;
        signal fifo_full_140095589934808: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140095589934808: core_fifo_inputs_t;
        signal outputs_full_140095589934808: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        

begin

    
        fifo_inputs_140095589890760(0) <= outputs_140095589890200(0);
        outputs_full_140095589890200(0) <= fifo_full_140095589890760(0);
        
        fifo_inputs_140095589890424(1) <= outputs_140095589890200(1);
        outputs_full_140095589890200(1) <= fifo_full_140095589890424(1);
        
        fifo_inputs_140095589890312(0) <= outputs_140095589890424(0);
        outputs_full_140095589890424(0) <= fifo_full_140095589890312(0);
        
        fifo_inputs_140095589890368(1) <= outputs_140095589890424(1);
        outputs_full_140095589890424(1) <= fifo_full_140095589890368(1);
        
        fifo_inputs_140095589890200(2) <= outputs_140095589890424(2);
        outputs_full_140095589890424(2) <= fifo_full_140095589890200(2);
        
        fifo_inputs_140095589890816(0) <= outputs_140095589890368(0);
        outputs_full_140095589890368(0) <= fifo_full_140095589890816(0);
        
        fifo_inputs_140095589890480(1) <= outputs_140095589890368(1);
        outputs_full_140095589890368(1) <= fifo_full_140095589890480(1);
        
        fifo_inputs_140095589890424(2) <= outputs_140095589890368(2);
        outputs_full_140095589890368(2) <= fifo_full_140095589890424(2);
        
        fifo_inputs_140095589890872(0) <= outputs_140095589890480(0);
        outputs_full_140095589890480(0) <= fifo_full_140095589890872(0);
        
        fifo_inputs_140095589890536(1) <= outputs_140095589890480(1);
        outputs_full_140095589890480(1) <= fifo_full_140095589890536(1);
        
        fifo_inputs_140095589890368(2) <= outputs_140095589890480(2);
        outputs_full_140095589890480(2) <= fifo_full_140095589890368(2);
        
        fifo_inputs_140095589890928(0) <= outputs_140095589890536(0);
        outputs_full_140095589890536(0) <= fifo_full_140095589890928(0);
        
        fifo_inputs_140095589890592(1) <= outputs_140095589890536(1);
        outputs_full_140095589890536(1) <= fifo_full_140095589890592(1);
        
        fifo_inputs_140095589890480(2) <= outputs_140095589890536(2);
        outputs_full_140095589890536(2) <= fifo_full_140095589890480(2);
        
        fifo_inputs_140095589890984(0) <= outputs_140095589890592(0);
        outputs_full_140095589890592(0) <= fifo_full_140095589890984(0);
        
        fifo_inputs_140095589890648(1) <= outputs_140095589890592(1);
        outputs_full_140095589890592(1) <= fifo_full_140095589890648(1);
        
        fifo_inputs_140095589890536(2) <= outputs_140095589890592(2);
        outputs_full_140095589890592(2) <= fifo_full_140095589890536(2);
        
        fifo_inputs_140095589891040(0) <= outputs_140095589890648(0);
        outputs_full_140095589890648(0) <= fifo_full_140095589891040(0);
        
        fifo_inputs_140095589890704(1) <= outputs_140095589890648(1);
        outputs_full_140095589890648(1) <= fifo_full_140095589890704(1);
        
        fifo_inputs_140095589890592(2) <= outputs_140095589890648(2);
        outputs_full_140095589890648(2) <= fifo_full_140095589890592(2);
        
        fifo_inputs_140095589891096(0) <= outputs_140095589890704(0);
        outputs_full_140095589890704(0) <= fifo_full_140095589891096(0);
        
        fifo_inputs_140095589890648(1) <= outputs_140095589890704(1);
        outputs_full_140095589890704(1) <= fifo_full_140095589890648(1);
        
        fifo_inputs_140095589891152(0) <= outputs_140095589890760(0);
        outputs_full_140095589890760(0) <= fifo_full_140095589891152(0);
        
        fifo_inputs_140095589890312(1) <= outputs_140095589890760(1);
        outputs_full_140095589890760(1) <= fifo_full_140095589890312(1);
        
        fifo_inputs_140095589890200(2) <= outputs_140095589890760(2);
        outputs_full_140095589890760(2) <= fifo_full_140095589890200(2);
        
        fifo_inputs_140095589891208(0) <= outputs_140095589890312(0);
        outputs_full_140095589890312(0) <= fifo_full_140095589891208(0);
        
        fifo_inputs_140095589890816(1) <= outputs_140095589890312(1);
        outputs_full_140095589890312(1) <= fifo_full_140095589890816(1);
        
        fifo_inputs_140095589890424(2) <= outputs_140095589890312(2);
        outputs_full_140095589890312(2) <= fifo_full_140095589890424(2);
        
        fifo_inputs_140095589890760(3) <= outputs_140095589890312(3);
        outputs_full_140095589890312(3) <= fifo_full_140095589890760(3);
        
        fifo_inputs_140095589891264(0) <= outputs_140095589890816(0);
        outputs_full_140095589890816(0) <= fifo_full_140095589891264(0);
        
        fifo_inputs_140095589890872(1) <= outputs_140095589890816(1);
        outputs_full_140095589890816(1) <= fifo_full_140095589890872(1);
        
        fifo_inputs_140095589890368(2) <= outputs_140095589890816(2);
        outputs_full_140095589890816(2) <= fifo_full_140095589890368(2);
        
        fifo_inputs_140095589890312(3) <= outputs_140095589890816(3);
        outputs_full_140095589890816(3) <= fifo_full_140095589890312(3);
        
        fifo_inputs_140095589891320(0) <= outputs_140095589890872(0);
        outputs_full_140095589890872(0) <= fifo_full_140095589891320(0);
        
        fifo_inputs_140095589890928(1) <= outputs_140095589890872(1);
        outputs_full_140095589890872(1) <= fifo_full_140095589890928(1);
        
        fifo_inputs_140095589890480(2) <= outputs_140095589890872(2);
        outputs_full_140095589890872(2) <= fifo_full_140095589890480(2);
        
        fifo_inputs_140095589890816(3) <= outputs_140095589890872(3);
        outputs_full_140095589890872(3) <= fifo_full_140095589890816(3);
        
        fifo_inputs_140095589891376(0) <= outputs_140095589890928(0);
        outputs_full_140095589890928(0) <= fifo_full_140095589891376(0);
        
        fifo_inputs_140095589890984(1) <= outputs_140095589890928(1);
        outputs_full_140095589890928(1) <= fifo_full_140095589890984(1);
        
        fifo_inputs_140095589890536(2) <= outputs_140095589890928(2);
        outputs_full_140095589890928(2) <= fifo_full_140095589890536(2);
        
        fifo_inputs_140095589890872(3) <= outputs_140095589890928(3);
        outputs_full_140095589890928(3) <= fifo_full_140095589890872(3);
        
        fifo_inputs_140095589891432(0) <= outputs_140095589890984(0);
        outputs_full_140095589890984(0) <= fifo_full_140095589891432(0);
        
        fifo_inputs_140095589891040(1) <= outputs_140095589890984(1);
        outputs_full_140095589890984(1) <= fifo_full_140095589891040(1);
        
        fifo_inputs_140095589890592(2) <= outputs_140095589890984(2);
        outputs_full_140095589890984(2) <= fifo_full_140095589890592(2);
        
        fifo_inputs_140095589890928(3) <= outputs_140095589890984(3);
        outputs_full_140095589890984(3) <= fifo_full_140095589890928(3);
        
        fifo_inputs_140095589891488(0) <= outputs_140095589891040(0);
        outputs_full_140095589891040(0) <= fifo_full_140095589891488(0);
        
        fifo_inputs_140095589891096(1) <= outputs_140095589891040(1);
        outputs_full_140095589891040(1) <= fifo_full_140095589891096(1);
        
        fifo_inputs_140095589890648(2) <= outputs_140095589891040(2);
        outputs_full_140095589891040(2) <= fifo_full_140095589890648(2);
        
        fifo_inputs_140095589890984(3) <= outputs_140095589891040(3);
        outputs_full_140095589891040(3) <= fifo_full_140095589890984(3);
        
        fifo_inputs_140095589891544(0) <= outputs_140095589891096(0);
        outputs_full_140095589891096(0) <= fifo_full_140095589891544(0);
        
        fifo_inputs_140095589890704(1) <= outputs_140095589891096(1);
        outputs_full_140095589891096(1) <= fifo_full_140095589890704(1);
        
        fifo_inputs_140095589891040(2) <= outputs_140095589891096(2);
        outputs_full_140095589891096(2) <= fifo_full_140095589891040(2);
        
        fifo_inputs_140095589891600(0) <= outputs_140095589891152(0);
        outputs_full_140095589891152(0) <= fifo_full_140095589891600(0);
        
        fifo_inputs_140095589891208(1) <= outputs_140095589891152(1);
        outputs_full_140095589891152(1) <= fifo_full_140095589891208(1);
        
        fifo_inputs_140095589890760(2) <= outputs_140095589891152(2);
        outputs_full_140095589891152(2) <= fifo_full_140095589890760(2);
        
        fifo_inputs_140095589891656(0) <= outputs_140095589891208(0);
        outputs_full_140095589891208(0) <= fifo_full_140095589891656(0);
        
        fifo_inputs_140095589891264(1) <= outputs_140095589891208(1);
        outputs_full_140095589891208(1) <= fifo_full_140095589891264(1);
        
        fifo_inputs_140095589890312(2) <= outputs_140095589891208(2);
        outputs_full_140095589891208(2) <= fifo_full_140095589890312(2);
        
        fifo_inputs_140095589891152(3) <= outputs_140095589891208(3);
        outputs_full_140095589891208(3) <= fifo_full_140095589891152(3);
        
        fifo_inputs_140095589891712(0) <= outputs_140095589891264(0);
        outputs_full_140095589891264(0) <= fifo_full_140095589891712(0);
        
        fifo_inputs_140095589891320(1) <= outputs_140095589891264(1);
        outputs_full_140095589891264(1) <= fifo_full_140095589891320(1);
        
        fifo_inputs_140095589890816(2) <= outputs_140095589891264(2);
        outputs_full_140095589891264(2) <= fifo_full_140095589890816(2);
        
        fifo_inputs_140095589891208(3) <= outputs_140095589891264(3);
        outputs_full_140095589891264(3) <= fifo_full_140095589891208(3);
        
        fifo_inputs_140095589891768(0) <= outputs_140095589891320(0);
        outputs_full_140095589891320(0) <= fifo_full_140095589891768(0);
        
        fifo_inputs_140095589891376(1) <= outputs_140095589891320(1);
        outputs_full_140095589891320(1) <= fifo_full_140095589891376(1);
        
        fifo_inputs_140095589890872(2) <= outputs_140095589891320(2);
        outputs_full_140095589891320(2) <= fifo_full_140095589890872(2);
        
        fifo_inputs_140095589891264(3) <= outputs_140095589891320(3);
        outputs_full_140095589891320(3) <= fifo_full_140095589891264(3);
        
        fifo_inputs_140095589891824(0) <= outputs_140095589891376(0);
        outputs_full_140095589891376(0) <= fifo_full_140095589891824(0);
        
        fifo_inputs_140095589891432(1) <= outputs_140095589891376(1);
        outputs_full_140095589891376(1) <= fifo_full_140095589891432(1);
        
        fifo_inputs_140095589890928(2) <= outputs_140095589891376(2);
        outputs_full_140095589891376(2) <= fifo_full_140095589890928(2);
        
        fifo_inputs_140095589891320(3) <= outputs_140095589891376(3);
        outputs_full_140095589891376(3) <= fifo_full_140095589891320(3);
        
        fifo_inputs_140095589891880(0) <= outputs_140095589891432(0);
        outputs_full_140095589891432(0) <= fifo_full_140095589891880(0);
        
        fifo_inputs_140095589891488(1) <= outputs_140095589891432(1);
        outputs_full_140095589891432(1) <= fifo_full_140095589891488(1);
        
        fifo_inputs_140095589890984(2) <= outputs_140095589891432(2);
        outputs_full_140095589891432(2) <= fifo_full_140095589890984(2);
        
        fifo_inputs_140095589891376(3) <= outputs_140095589891432(3);
        outputs_full_140095589891432(3) <= fifo_full_140095589891376(3);
        
        fifo_inputs_140095589891936(0) <= outputs_140095589891488(0);
        outputs_full_140095589891488(0) <= fifo_full_140095589891936(0);
        
        fifo_inputs_140095589891544(1) <= outputs_140095589891488(1);
        outputs_full_140095589891488(1) <= fifo_full_140095589891544(1);
        
        fifo_inputs_140095589891040(2) <= outputs_140095589891488(2);
        outputs_full_140095589891488(2) <= fifo_full_140095589891040(2);
        
        fifo_inputs_140095589891432(3) <= outputs_140095589891488(3);
        outputs_full_140095589891488(3) <= fifo_full_140095589891432(3);
        
        fifo_inputs_140095589891992(0) <= outputs_140095589891544(0);
        outputs_full_140095589891544(0) <= fifo_full_140095589891992(0);
        
        fifo_inputs_140095589891096(1) <= outputs_140095589891544(1);
        outputs_full_140095589891544(1) <= fifo_full_140095589891096(1);
        
        fifo_inputs_140095589891488(2) <= outputs_140095589891544(2);
        outputs_full_140095589891544(2) <= fifo_full_140095589891488(2);
        
        fifo_inputs_140095589892048(0) <= outputs_140095589891600(0);
        outputs_full_140095589891600(0) <= fifo_full_140095589892048(0);
        
        fifo_inputs_140095589891656(1) <= outputs_140095589891600(1);
        outputs_full_140095589891600(1) <= fifo_full_140095589891656(1);
        
        fifo_inputs_140095589891152(2) <= outputs_140095589891600(2);
        outputs_full_140095589891600(2) <= fifo_full_140095589891152(2);
        
        fifo_inputs_140095589933128(0) <= outputs_140095589891656(0);
        outputs_full_140095589891656(0) <= fifo_full_140095589933128(0);
        
        fifo_inputs_140095589891712(1) <= outputs_140095589891656(1);
        outputs_full_140095589891656(1) <= fifo_full_140095589891712(1);
        
        fifo_inputs_140095589891208(2) <= outputs_140095589891656(2);
        outputs_full_140095589891656(2) <= fifo_full_140095589891208(2);
        
        fifo_inputs_140095589891600(3) <= outputs_140095589891656(3);
        outputs_full_140095589891656(3) <= fifo_full_140095589891600(3);
        
        fifo_inputs_140095589933184(0) <= outputs_140095589891712(0);
        outputs_full_140095589891712(0) <= fifo_full_140095589933184(0);
        
        fifo_inputs_140095589891768(1) <= outputs_140095589891712(1);
        outputs_full_140095589891712(1) <= fifo_full_140095589891768(1);
        
        fifo_inputs_140095589891264(2) <= outputs_140095589891712(2);
        outputs_full_140095589891712(2) <= fifo_full_140095589891264(2);
        
        fifo_inputs_140095589891656(3) <= outputs_140095589891712(3);
        outputs_full_140095589891712(3) <= fifo_full_140095589891656(3);
        
        fifo_inputs_140095589933240(0) <= outputs_140095589891768(0);
        outputs_full_140095589891768(0) <= fifo_full_140095589933240(0);
        
        fifo_inputs_140095589891824(1) <= outputs_140095589891768(1);
        outputs_full_140095589891768(1) <= fifo_full_140095589891824(1);
        
        fifo_inputs_140095589891320(2) <= outputs_140095589891768(2);
        outputs_full_140095589891768(2) <= fifo_full_140095589891320(2);
        
        fifo_inputs_140095589891712(3) <= outputs_140095589891768(3);
        outputs_full_140095589891768(3) <= fifo_full_140095589891712(3);
        
        fifo_inputs_140095589933296(0) <= outputs_140095589891824(0);
        outputs_full_140095589891824(0) <= fifo_full_140095589933296(0);
        
        fifo_inputs_140095589891880(1) <= outputs_140095589891824(1);
        outputs_full_140095589891824(1) <= fifo_full_140095589891880(1);
        
        fifo_inputs_140095589891376(2) <= outputs_140095589891824(2);
        outputs_full_140095589891824(2) <= fifo_full_140095589891376(2);
        
        fifo_inputs_140095589891768(3) <= outputs_140095589891824(3);
        outputs_full_140095589891824(3) <= fifo_full_140095589891768(3);
        
        fifo_inputs_140095589933352(0) <= outputs_140095589891880(0);
        outputs_full_140095589891880(0) <= fifo_full_140095589933352(0);
        
        fifo_inputs_140095589891936(1) <= outputs_140095589891880(1);
        outputs_full_140095589891880(1) <= fifo_full_140095589891936(1);
        
        fifo_inputs_140095589891432(2) <= outputs_140095589891880(2);
        outputs_full_140095589891880(2) <= fifo_full_140095589891432(2);
        
        fifo_inputs_140095589891824(3) <= outputs_140095589891880(3);
        outputs_full_140095589891880(3) <= fifo_full_140095589891824(3);
        
        fifo_inputs_140095589933408(0) <= outputs_140095589891936(0);
        outputs_full_140095589891936(0) <= fifo_full_140095589933408(0);
        
        fifo_inputs_140095589891992(1) <= outputs_140095589891936(1);
        outputs_full_140095589891936(1) <= fifo_full_140095589891992(1);
        
        fifo_inputs_140095589891488(2) <= outputs_140095589891936(2);
        outputs_full_140095589891936(2) <= fifo_full_140095589891488(2);
        
        fifo_inputs_140095589891880(3) <= outputs_140095589891936(3);
        outputs_full_140095589891936(3) <= fifo_full_140095589891880(3);
        
        fifo_inputs_140095589933464(0) <= outputs_140095589891992(0);
        outputs_full_140095589891992(0) <= fifo_full_140095589933464(0);
        
        fifo_inputs_140095589891544(1) <= outputs_140095589891992(1);
        outputs_full_140095589891992(1) <= fifo_full_140095589891544(1);
        
        fifo_inputs_140095589891936(2) <= outputs_140095589891992(2);
        outputs_full_140095589891992(2) <= fifo_full_140095589891936(2);
        
        fifo_inputs_140095589933520(0) <= outputs_140095589892048(0);
        outputs_full_140095589892048(0) <= fifo_full_140095589933520(0);
        
        fifo_inputs_140095589933128(1) <= outputs_140095589892048(1);
        outputs_full_140095589892048(1) <= fifo_full_140095589933128(1);
        
        fifo_inputs_140095589891600(2) <= outputs_140095589892048(2);
        outputs_full_140095589892048(2) <= fifo_full_140095589891600(2);
        
        fifo_inputs_140095589933576(0) <= outputs_140095589933128(0);
        outputs_full_140095589933128(0) <= fifo_full_140095589933576(0);
        
        fifo_inputs_140095589933184(1) <= outputs_140095589933128(1);
        outputs_full_140095589933128(1) <= fifo_full_140095589933184(1);
        
        fifo_inputs_140095589891656(2) <= outputs_140095589933128(2);
        outputs_full_140095589933128(2) <= fifo_full_140095589891656(2);
        
        fifo_inputs_140095589892048(3) <= outputs_140095589933128(3);
        outputs_full_140095589933128(3) <= fifo_full_140095589892048(3);
        
        fifo_inputs_140095589933632(0) <= outputs_140095589933184(0);
        outputs_full_140095589933184(0) <= fifo_full_140095589933632(0);
        
        fifo_inputs_140095589933240(1) <= outputs_140095589933184(1);
        outputs_full_140095589933184(1) <= fifo_full_140095589933240(1);
        
        fifo_inputs_140095589891712(2) <= outputs_140095589933184(2);
        outputs_full_140095589933184(2) <= fifo_full_140095589891712(2);
        
        fifo_inputs_140095589933128(3) <= outputs_140095589933184(3);
        outputs_full_140095589933184(3) <= fifo_full_140095589933128(3);
        
        fifo_inputs_140095589933688(0) <= outputs_140095589933240(0);
        outputs_full_140095589933240(0) <= fifo_full_140095589933688(0);
        
        fifo_inputs_140095589933296(1) <= outputs_140095589933240(1);
        outputs_full_140095589933240(1) <= fifo_full_140095589933296(1);
        
        fifo_inputs_140095589891768(2) <= outputs_140095589933240(2);
        outputs_full_140095589933240(2) <= fifo_full_140095589891768(2);
        
        fifo_inputs_140095589933184(3) <= outputs_140095589933240(3);
        outputs_full_140095589933240(3) <= fifo_full_140095589933184(3);
        
        fifo_inputs_140095589933744(0) <= outputs_140095589933296(0);
        outputs_full_140095589933296(0) <= fifo_full_140095589933744(0);
        
        fifo_inputs_140095589933352(1) <= outputs_140095589933296(1);
        outputs_full_140095589933296(1) <= fifo_full_140095589933352(1);
        
        fifo_inputs_140095589891824(2) <= outputs_140095589933296(2);
        outputs_full_140095589933296(2) <= fifo_full_140095589891824(2);
        
        fifo_inputs_140095589933240(3) <= outputs_140095589933296(3);
        outputs_full_140095589933296(3) <= fifo_full_140095589933240(3);
        
        fifo_inputs_140095589933800(0) <= outputs_140095589933352(0);
        outputs_full_140095589933352(0) <= fifo_full_140095589933800(0);
        
        fifo_inputs_140095589933408(1) <= outputs_140095589933352(1);
        outputs_full_140095589933352(1) <= fifo_full_140095589933408(1);
        
        fifo_inputs_140095589891880(2) <= outputs_140095589933352(2);
        outputs_full_140095589933352(2) <= fifo_full_140095589891880(2);
        
        fifo_inputs_140095589933296(3) <= outputs_140095589933352(3);
        outputs_full_140095589933352(3) <= fifo_full_140095589933296(3);
        
        fifo_inputs_140095589933856(0) <= outputs_140095589933408(0);
        outputs_full_140095589933408(0) <= fifo_full_140095589933856(0);
        
        fifo_inputs_140095589933464(1) <= outputs_140095589933408(1);
        outputs_full_140095589933408(1) <= fifo_full_140095589933464(1);
        
        fifo_inputs_140095589891936(2) <= outputs_140095589933408(2);
        outputs_full_140095589933408(2) <= fifo_full_140095589891936(2);
        
        fifo_inputs_140095589933352(3) <= outputs_140095589933408(3);
        outputs_full_140095589933408(3) <= fifo_full_140095589933352(3);
        
        fifo_inputs_140095589933912(0) <= outputs_140095589933464(0);
        outputs_full_140095589933464(0) <= fifo_full_140095589933912(0);
        
        fifo_inputs_140095589891992(1) <= outputs_140095589933464(1);
        outputs_full_140095589933464(1) <= fifo_full_140095589891992(1);
        
        fifo_inputs_140095589933408(2) <= outputs_140095589933464(2);
        outputs_full_140095589933464(2) <= fifo_full_140095589933408(2);
        
        fifo_inputs_140095589933968(0) <= outputs_140095589933520(0);
        outputs_full_140095589933520(0) <= fifo_full_140095589933968(0);
        
        fifo_inputs_140095589933576(1) <= outputs_140095589933520(1);
        outputs_full_140095589933520(1) <= fifo_full_140095589933576(1);
        
        fifo_inputs_140095589892048(2) <= outputs_140095589933520(2);
        outputs_full_140095589933520(2) <= fifo_full_140095589892048(2);
        
        fifo_inputs_140095589934024(0) <= outputs_140095589933576(0);
        outputs_full_140095589933576(0) <= fifo_full_140095589934024(0);
        
        fifo_inputs_140095589933632(1) <= outputs_140095589933576(1);
        outputs_full_140095589933576(1) <= fifo_full_140095589933632(1);
        
        fifo_inputs_140095589933128(2) <= outputs_140095589933576(2);
        outputs_full_140095589933576(2) <= fifo_full_140095589933128(2);
        
        fifo_inputs_140095589933520(3) <= outputs_140095589933576(3);
        outputs_full_140095589933576(3) <= fifo_full_140095589933520(3);
        
        fifo_inputs_140095589934080(0) <= outputs_140095589933632(0);
        outputs_full_140095589933632(0) <= fifo_full_140095589934080(0);
        
        fifo_inputs_140095589933688(1) <= outputs_140095589933632(1);
        outputs_full_140095589933632(1) <= fifo_full_140095589933688(1);
        
        fifo_inputs_140095589933184(2) <= outputs_140095589933632(2);
        outputs_full_140095589933632(2) <= fifo_full_140095589933184(2);
        
        fifo_inputs_140095589933576(3) <= outputs_140095589933632(3);
        outputs_full_140095589933632(3) <= fifo_full_140095589933576(3);
        
        fifo_inputs_140095589934136(0) <= outputs_140095589933688(0);
        outputs_full_140095589933688(0) <= fifo_full_140095589934136(0);
        
        fifo_inputs_140095589933744(1) <= outputs_140095589933688(1);
        outputs_full_140095589933688(1) <= fifo_full_140095589933744(1);
        
        fifo_inputs_140095589933240(2) <= outputs_140095589933688(2);
        outputs_full_140095589933688(2) <= fifo_full_140095589933240(2);
        
        fifo_inputs_140095589933632(3) <= outputs_140095589933688(3);
        outputs_full_140095589933688(3) <= fifo_full_140095589933632(3);
        
        fifo_inputs_140095589934192(0) <= outputs_140095589933744(0);
        outputs_full_140095589933744(0) <= fifo_full_140095589934192(0);
        
        fifo_inputs_140095589933800(1) <= outputs_140095589933744(1);
        outputs_full_140095589933744(1) <= fifo_full_140095589933800(1);
        
        fifo_inputs_140095589933296(2) <= outputs_140095589933744(2);
        outputs_full_140095589933744(2) <= fifo_full_140095589933296(2);
        
        fifo_inputs_140095589933688(3) <= outputs_140095589933744(3);
        outputs_full_140095589933744(3) <= fifo_full_140095589933688(3);
        
        fifo_inputs_140095589934248(0) <= outputs_140095589933800(0);
        outputs_full_140095589933800(0) <= fifo_full_140095589934248(0);
        
        fifo_inputs_140095589933856(1) <= outputs_140095589933800(1);
        outputs_full_140095589933800(1) <= fifo_full_140095589933856(1);
        
        fifo_inputs_140095589933352(2) <= outputs_140095589933800(2);
        outputs_full_140095589933800(2) <= fifo_full_140095589933352(2);
        
        fifo_inputs_140095589933744(3) <= outputs_140095589933800(3);
        outputs_full_140095589933800(3) <= fifo_full_140095589933744(3);
        
        fifo_inputs_140095589934304(0) <= outputs_140095589933856(0);
        outputs_full_140095589933856(0) <= fifo_full_140095589934304(0);
        
        fifo_inputs_140095589933912(1) <= outputs_140095589933856(1);
        outputs_full_140095589933856(1) <= fifo_full_140095589933912(1);
        
        fifo_inputs_140095589933408(2) <= outputs_140095589933856(2);
        outputs_full_140095589933856(2) <= fifo_full_140095589933408(2);
        
        fifo_inputs_140095589933800(3) <= outputs_140095589933856(3);
        outputs_full_140095589933856(3) <= fifo_full_140095589933800(3);
        
        fifo_inputs_140095589934360(0) <= outputs_140095589933912(0);
        outputs_full_140095589933912(0) <= fifo_full_140095589934360(0);
        
        fifo_inputs_140095589933464(1) <= outputs_140095589933912(1);
        outputs_full_140095589933912(1) <= fifo_full_140095589933464(1);
        
        fifo_inputs_140095589933856(2) <= outputs_140095589933912(2);
        outputs_full_140095589933912(2) <= fifo_full_140095589933856(2);
        
        fifo_inputs_140095589934416(0) <= outputs_140095589933968(0);
        outputs_full_140095589933968(0) <= fifo_full_140095589934416(0);
        
        fifo_inputs_140095589934024(1) <= outputs_140095589933968(1);
        outputs_full_140095589933968(1) <= fifo_full_140095589934024(1);
        
        fifo_inputs_140095589933520(2) <= outputs_140095589933968(2);
        outputs_full_140095589933968(2) <= fifo_full_140095589933520(2);
        
        fifo_inputs_140095589934472(0) <= outputs_140095589934024(0);
        outputs_full_140095589934024(0) <= fifo_full_140095589934472(0);
        
        fifo_inputs_140095589934080(1) <= outputs_140095589934024(1);
        outputs_full_140095589934024(1) <= fifo_full_140095589934080(1);
        
        fifo_inputs_140095589933576(2) <= outputs_140095589934024(2);
        outputs_full_140095589934024(2) <= fifo_full_140095589933576(2);
        
        fifo_inputs_140095589933968(3) <= outputs_140095589934024(3);
        outputs_full_140095589934024(3) <= fifo_full_140095589933968(3);
        
        fifo_inputs_140095589934528(0) <= outputs_140095589934080(0);
        outputs_full_140095589934080(0) <= fifo_full_140095589934528(0);
        
        fifo_inputs_140095589934136(1) <= outputs_140095589934080(1);
        outputs_full_140095589934080(1) <= fifo_full_140095589934136(1);
        
        fifo_inputs_140095589933632(2) <= outputs_140095589934080(2);
        outputs_full_140095589934080(2) <= fifo_full_140095589933632(2);
        
        fifo_inputs_140095589934024(3) <= outputs_140095589934080(3);
        outputs_full_140095589934080(3) <= fifo_full_140095589934024(3);
        
        fifo_inputs_140095589934584(0) <= outputs_140095589934136(0);
        outputs_full_140095589934136(0) <= fifo_full_140095589934584(0);
        
        fifo_inputs_140095589934192(1) <= outputs_140095589934136(1);
        outputs_full_140095589934136(1) <= fifo_full_140095589934192(1);
        
        fifo_inputs_140095589933688(2) <= outputs_140095589934136(2);
        outputs_full_140095589934136(2) <= fifo_full_140095589933688(2);
        
        fifo_inputs_140095589934080(3) <= outputs_140095589934136(3);
        outputs_full_140095589934136(3) <= fifo_full_140095589934080(3);
        
        fifo_inputs_140095589934640(0) <= outputs_140095589934192(0);
        outputs_full_140095589934192(0) <= fifo_full_140095589934640(0);
        
        fifo_inputs_140095589934248(1) <= outputs_140095589934192(1);
        outputs_full_140095589934192(1) <= fifo_full_140095589934248(1);
        
        fifo_inputs_140095589933744(2) <= outputs_140095589934192(2);
        outputs_full_140095589934192(2) <= fifo_full_140095589933744(2);
        
        fifo_inputs_140095589934136(3) <= outputs_140095589934192(3);
        outputs_full_140095589934192(3) <= fifo_full_140095589934136(3);
        
        fifo_inputs_140095589934696(0) <= outputs_140095589934248(0);
        outputs_full_140095589934248(0) <= fifo_full_140095589934696(0);
        
        fifo_inputs_140095589934304(1) <= outputs_140095589934248(1);
        outputs_full_140095589934248(1) <= fifo_full_140095589934304(1);
        
        fifo_inputs_140095589933800(2) <= outputs_140095589934248(2);
        outputs_full_140095589934248(2) <= fifo_full_140095589933800(2);
        
        fifo_inputs_140095589934192(3) <= outputs_140095589934248(3);
        outputs_full_140095589934248(3) <= fifo_full_140095589934192(3);
        
        fifo_inputs_140095589934752(0) <= outputs_140095589934304(0);
        outputs_full_140095589934304(0) <= fifo_full_140095589934752(0);
        
        fifo_inputs_140095589934360(1) <= outputs_140095589934304(1);
        outputs_full_140095589934304(1) <= fifo_full_140095589934360(1);
        
        fifo_inputs_140095589933856(2) <= outputs_140095589934304(2);
        outputs_full_140095589934304(2) <= fifo_full_140095589933856(2);
        
        fifo_inputs_140095589934248(3) <= outputs_140095589934304(3);
        outputs_full_140095589934304(3) <= fifo_full_140095589934248(3);
        
        fifo_inputs_140095589934808(0) <= outputs_140095589934360(0);
        outputs_full_140095589934360(0) <= fifo_full_140095589934808(0);
        
        fifo_inputs_140095589933912(1) <= outputs_140095589934360(1);
        outputs_full_140095589934360(1) <= fifo_full_140095589933912(1);
        
        fifo_inputs_140095589934304(2) <= outputs_140095589934360(2);
        outputs_full_140095589934360(2) <= fifo_full_140095589934304(2);
        
        fifo_inputs_140095589934472(0) <= outputs_140095589934416(0);
        outputs_full_140095589934416(0) <= fifo_full_140095589934472(0);
        
        fifo_inputs_140095589933968(1) <= outputs_140095589934416(1);
        outputs_full_140095589934416(1) <= fifo_full_140095589933968(1);
        
        fifo_inputs_140095589934528(0) <= outputs_140095589934472(0);
        outputs_full_140095589934472(0) <= fifo_full_140095589934528(0);
        
        fifo_inputs_140095589934024(1) <= outputs_140095589934472(1);
        outputs_full_140095589934472(1) <= fifo_full_140095589934024(1);
        
        fifo_inputs_140095589934416(2) <= outputs_140095589934472(2);
        outputs_full_140095589934472(2) <= fifo_full_140095589934416(2);
        
        fifo_inputs_140095589934584(0) <= outputs_140095589934528(0);
        outputs_full_140095589934528(0) <= fifo_full_140095589934584(0);
        
        fifo_inputs_140095589934080(1) <= outputs_140095589934528(1);
        outputs_full_140095589934528(1) <= fifo_full_140095589934080(1);
        
        fifo_inputs_140095589934472(2) <= outputs_140095589934528(2);
        outputs_full_140095589934528(2) <= fifo_full_140095589934472(2);
        
        fifo_inputs_140095589934640(0) <= outputs_140095589934584(0);
        outputs_full_140095589934584(0) <= fifo_full_140095589934640(0);
        
        fifo_inputs_140095589934136(1) <= outputs_140095589934584(1);
        outputs_full_140095589934584(1) <= fifo_full_140095589934136(1);
        
        fifo_inputs_140095589934528(2) <= outputs_140095589934584(2);
        outputs_full_140095589934584(2) <= fifo_full_140095589934528(2);
        
        fifo_inputs_140095589934696(0) <= outputs_140095589934640(0);
        outputs_full_140095589934640(0) <= fifo_full_140095589934696(0);
        
        fifo_inputs_140095589934192(1) <= outputs_140095589934640(1);
        outputs_full_140095589934640(1) <= fifo_full_140095589934192(1);
        
        fifo_inputs_140095589934584(2) <= outputs_140095589934640(2);
        outputs_full_140095589934640(2) <= fifo_full_140095589934584(2);
        
        fifo_inputs_140095589934752(0) <= outputs_140095589934696(0);
        outputs_full_140095589934696(0) <= fifo_full_140095589934752(0);
        
        fifo_inputs_140095589934248(1) <= outputs_140095589934696(1);
        outputs_full_140095589934696(1) <= fifo_full_140095589934248(1);
        
        fifo_inputs_140095589934640(2) <= outputs_140095589934696(2);
        outputs_full_140095589934696(2) <= fifo_full_140095589934640(2);
        
        fifo_inputs_140095589934808(0) <= outputs_140095589934752(0);
        outputs_full_140095589934752(0) <= fifo_full_140095589934808(0);
        
        fifo_inputs_140095589934304(1) <= outputs_140095589934752(1);
        outputs_full_140095589934752(1) <= fifo_full_140095589934304(1);
        
        fifo_inputs_140095589934696(2) <= outputs_140095589934752(2);
        outputs_full_140095589934752(2) <= fifo_full_140095589934696(2);
        
        fifo_inputs_140095589934360(0) <= outputs_140095589934808(0);
        outputs_full_140095589934808(0) <= fifo_full_140095589934360(0);
        
        fifo_inputs_140095589934752(1) <= outputs_140095589934808(1);
        outputs_full_140095589934808(1) <= fifo_full_140095589934752(1);
        

    
        core_inst_140095589890200: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589890200,
            fifo_full => fifo_full_140095589890200,
            outputs => outputs_140095589890200,
            outputs_full => outputs_full_140095589890200
        );
        
        core_inst_140095589890424: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589890424,
            fifo_full => fifo_full_140095589890424,
            outputs => outputs_140095589890424,
            outputs_full => outputs_full_140095589890424
        );
        
        core_inst_140095589890368: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589890368,
            fifo_full => fifo_full_140095589890368,
            outputs => outputs_140095589890368,
            outputs_full => outputs_full_140095589890368
        );
        
        core_inst_140095589890480: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589890480,
            fifo_full => fifo_full_140095589890480,
            outputs => outputs_140095589890480,
            outputs_full => outputs_full_140095589890480
        );
        
        core_inst_140095589890536: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589890536,
            fifo_full => fifo_full_140095589890536,
            outputs => outputs_140095589890536,
            outputs_full => outputs_full_140095589890536
        );
        
        core_inst_140095589890592: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589890592,
            fifo_full => fifo_full_140095589890592,
            outputs => outputs_140095589890592,
            outputs_full => outputs_full_140095589890592
        );
        
        core_inst_140095589890648: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589890648,
            fifo_full => fifo_full_140095589890648,
            outputs => outputs_140095589890648,
            outputs_full => outputs_full_140095589890648
        );
        
        core_inst_140095589890704: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589890704,
            fifo_full => fifo_full_140095589890704,
            outputs => outputs_140095589890704,
            outputs_full => outputs_full_140095589890704
        );
        
        core_inst_140095589890760: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589890760,
            fifo_full => fifo_full_140095589890760,
            outputs => outputs_140095589890760,
            outputs_full => outputs_full_140095589890760
        );
        
        core_inst_140095589890312: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589890312,
            fifo_full => fifo_full_140095589890312,
            outputs => outputs_140095589890312,
            outputs_full => outputs_full_140095589890312
        );
        
        core_inst_140095589890816: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589890816,
            fifo_full => fifo_full_140095589890816,
            outputs => outputs_140095589890816,
            outputs_full => outputs_full_140095589890816
        );
        
        core_inst_140095589890872: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589890872,
            fifo_full => fifo_full_140095589890872,
            outputs => outputs_140095589890872,
            outputs_full => outputs_full_140095589890872
        );
        
        core_inst_140095589890928: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589890928,
            fifo_full => fifo_full_140095589890928,
            outputs => outputs_140095589890928,
            outputs_full => outputs_full_140095589890928
        );
        
        core_inst_140095589890984: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589890984,
            fifo_full => fifo_full_140095589890984,
            outputs => outputs_140095589890984,
            outputs_full => outputs_full_140095589890984
        );
        
        core_inst_140095589891040: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589891040,
            fifo_full => fifo_full_140095589891040,
            outputs => outputs_140095589891040,
            outputs_full => outputs_full_140095589891040
        );
        
        core_inst_140095589891096: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589891096,
            fifo_full => fifo_full_140095589891096,
            outputs => outputs_140095589891096,
            outputs_full => outputs_full_140095589891096
        );
        
        core_inst_140095589891152: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589891152,
            fifo_full => fifo_full_140095589891152,
            outputs => outputs_140095589891152,
            outputs_full => outputs_full_140095589891152
        );
        
        core_inst_140095589891208: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589891208,
            fifo_full => fifo_full_140095589891208,
            outputs => outputs_140095589891208,
            outputs_full => outputs_full_140095589891208
        );
        
        core_inst_140095589891264: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589891264,
            fifo_full => fifo_full_140095589891264,
            outputs => outputs_140095589891264,
            outputs_full => outputs_full_140095589891264
        );
        
        core_inst_140095589891320: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589891320,
            fifo_full => fifo_full_140095589891320,
            outputs => outputs_140095589891320,
            outputs_full => outputs_full_140095589891320
        );
        
        core_inst_140095589891376: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589891376,
            fifo_full => fifo_full_140095589891376,
            outputs => outputs_140095589891376,
            outputs_full => outputs_full_140095589891376
        );
        
        core_inst_140095589891432: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589891432,
            fifo_full => fifo_full_140095589891432,
            outputs => outputs_140095589891432,
            outputs_full => outputs_full_140095589891432
        );
        
        core_inst_140095589891488: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589891488,
            fifo_full => fifo_full_140095589891488,
            outputs => outputs_140095589891488,
            outputs_full => outputs_full_140095589891488
        );
        
        core_inst_140095589891544: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589891544,
            fifo_full => fifo_full_140095589891544,
            outputs => outputs_140095589891544,
            outputs_full => outputs_full_140095589891544
        );
        
        core_inst_140095589891600: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589891600,
            fifo_full => fifo_full_140095589891600,
            outputs => outputs_140095589891600,
            outputs_full => outputs_full_140095589891600
        );
        
        core_inst_140095589891656: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589891656,
            fifo_full => fifo_full_140095589891656,
            outputs => outputs_140095589891656,
            outputs_full => outputs_full_140095589891656
        );
        
        core_inst_140095589891712: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589891712,
            fifo_full => fifo_full_140095589891712,
            outputs => outputs_140095589891712,
            outputs_full => outputs_full_140095589891712
        );
        
        core_inst_140095589891768: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589891768,
            fifo_full => fifo_full_140095589891768,
            outputs => outputs_140095589891768,
            outputs_full => outputs_full_140095589891768
        );
        
        core_inst_140095589891824: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589891824,
            fifo_full => fifo_full_140095589891824,
            outputs => outputs_140095589891824,
            outputs_full => outputs_full_140095589891824
        );
        
        core_inst_140095589891880: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589891880,
            fifo_full => fifo_full_140095589891880,
            outputs => outputs_140095589891880,
            outputs_full => outputs_full_140095589891880
        );
        
        core_inst_140095589891936: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589891936,
            fifo_full => fifo_full_140095589891936,
            outputs => outputs_140095589891936,
            outputs_full => outputs_full_140095589891936
        );
        
        core_inst_140095589891992: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589891992,
            fifo_full => fifo_full_140095589891992,
            outputs => outputs_140095589891992,
            outputs_full => outputs_full_140095589891992
        );
        
        core_inst_140095589892048: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589892048,
            fifo_full => fifo_full_140095589892048,
            outputs => outputs_140095589892048,
            outputs_full => outputs_full_140095589892048
        );
        
        core_inst_140095589933128: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589933128,
            fifo_full => fifo_full_140095589933128,
            outputs => outputs_140095589933128,
            outputs_full => outputs_full_140095589933128
        );
        
        core_inst_140095589933184: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589933184,
            fifo_full => fifo_full_140095589933184,
            outputs => outputs_140095589933184,
            outputs_full => outputs_full_140095589933184
        );
        
        core_inst_140095589933240: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589933240,
            fifo_full => fifo_full_140095589933240,
            outputs => outputs_140095589933240,
            outputs_full => outputs_full_140095589933240
        );
        
        core_inst_140095589933296: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589933296,
            fifo_full => fifo_full_140095589933296,
            outputs => outputs_140095589933296,
            outputs_full => outputs_full_140095589933296
        );
        
        core_inst_140095589933352: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589933352,
            fifo_full => fifo_full_140095589933352,
            outputs => outputs_140095589933352,
            outputs_full => outputs_full_140095589933352
        );
        
        core_inst_140095589933408: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589933408,
            fifo_full => fifo_full_140095589933408,
            outputs => outputs_140095589933408,
            outputs_full => outputs_full_140095589933408
        );
        
        core_inst_140095589933464: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589933464,
            fifo_full => fifo_full_140095589933464,
            outputs => outputs_140095589933464,
            outputs_full => outputs_full_140095589933464
        );
        
        core_inst_140095589933520: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589933520,
            fifo_full => fifo_full_140095589933520,
            outputs => outputs_140095589933520,
            outputs_full => outputs_full_140095589933520
        );
        
        core_inst_140095589933576: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589933576,
            fifo_full => fifo_full_140095589933576,
            outputs => outputs_140095589933576,
            outputs_full => outputs_full_140095589933576
        );
        
        core_inst_140095589933632: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589933632,
            fifo_full => fifo_full_140095589933632,
            outputs => outputs_140095589933632,
            outputs_full => outputs_full_140095589933632
        );
        
        core_inst_140095589933688: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589933688,
            fifo_full => fifo_full_140095589933688,
            outputs => outputs_140095589933688,
            outputs_full => outputs_full_140095589933688
        );
        
        core_inst_140095589933744: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589933744,
            fifo_full => fifo_full_140095589933744,
            outputs => outputs_140095589933744,
            outputs_full => outputs_full_140095589933744
        );
        
        core_inst_140095589933800: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589933800,
            fifo_full => fifo_full_140095589933800,
            outputs => outputs_140095589933800,
            outputs_full => outputs_full_140095589933800
        );
        
        core_inst_140095589933856: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589933856,
            fifo_full => fifo_full_140095589933856,
            outputs => outputs_140095589933856,
            outputs_full => outputs_full_140095589933856
        );
        
        core_inst_140095589933912: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589933912,
            fifo_full => fifo_full_140095589933912,
            outputs => outputs_140095589933912,
            outputs_full => outputs_full_140095589933912
        );
        
        core_inst_140095589933968: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589933968,
            fifo_full => fifo_full_140095589933968,
            outputs => outputs_140095589933968,
            outputs_full => outputs_full_140095589933968
        );
        
        core_inst_140095589934024: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589934024,
            fifo_full => fifo_full_140095589934024,
            outputs => outputs_140095589934024,
            outputs_full => outputs_full_140095589934024
        );
        
        core_inst_140095589934080: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589934080,
            fifo_full => fifo_full_140095589934080,
            outputs => outputs_140095589934080,
            outputs_full => outputs_full_140095589934080
        );
        
        core_inst_140095589934136: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589934136,
            fifo_full => fifo_full_140095589934136,
            outputs => outputs_140095589934136,
            outputs_full => outputs_full_140095589934136
        );
        
        core_inst_140095589934192: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589934192,
            fifo_full => fifo_full_140095589934192,
            outputs => outputs_140095589934192,
            outputs_full => outputs_full_140095589934192
        );
        
        core_inst_140095589934248: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589934248,
            fifo_full => fifo_full_140095589934248,
            outputs => outputs_140095589934248,
            outputs_full => outputs_full_140095589934248
        );
        
        core_inst_140095589934304: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589934304,
            fifo_full => fifo_full_140095589934304,
            outputs => outputs_140095589934304,
            outputs_full => outputs_full_140095589934304
        );
        
        core_inst_140095589934360: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589934360,
            fifo_full => fifo_full_140095589934360,
            outputs => outputs_140095589934360,
            outputs_full => outputs_full_140095589934360
        );
        
        core_inst_140095589934416: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589934416,
            fifo_full => fifo_full_140095589934416,
            outputs => outputs_140095589934416,
            outputs_full => outputs_full_140095589934416
        );
        
        core_inst_140095589934472: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589934472,
            fifo_full => fifo_full_140095589934472,
            outputs => outputs_140095589934472,
            outputs_full => outputs_full_140095589934472
        );
        
        core_inst_140095589934528: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589934528,
            fifo_full => fifo_full_140095589934528,
            outputs => outputs_140095589934528,
            outputs_full => outputs_full_140095589934528
        );
        
        core_inst_140095589934584: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589934584,
            fifo_full => fifo_full_140095589934584,
            outputs => outputs_140095589934584,
            outputs_full => outputs_full_140095589934584
        );
        
        core_inst_140095589934640: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589934640,
            fifo_full => fifo_full_140095589934640,
            outputs => outputs_140095589934640,
            outputs_full => outputs_full_140095589934640
        );
        
        core_inst_140095589934696: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589934696,
            fifo_full => fifo_full_140095589934696,
            outputs => outputs_140095589934696,
            outputs_full => outputs_full_140095589934696
        );
        
        core_inst_140095589934752: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589934752,
            fifo_full => fifo_full_140095589934752,
            outputs => outputs_140095589934752,
            outputs_full => outputs_full_140095589934752
        );
        
        core_inst_140095589934808: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140095589934808,
            fifo_full => fifo_full_140095589934808,
            outputs => outputs_140095589934808,
            outputs_full => outputs_full_140095589934808
        );
        

end behav;

