
library ieee;
use ieee.std_logic_1164.all;
use work.core_config.all;
use work.all;

entity Chain800 is
    port (
        clk: in std_logic;
        clk_en: in std_logic;
        reset: in std_logic;
        addr: in ram_addr;
        data: in word;
        we: in std_logic;
        fifo_inputs: in core_fifo_inputs_t;
        fifo_full: out std_logic_vector(0 to NUM_CORE_FIFOS-1);
        outputs: out core_fifo_inputs_t;
        outputs_full: in std_logic_vector(0 to NUM_CORE_FIFOS-1)
    );
end Chain800;

architecture behav of Chain800 is

    
        signal fifo_inputs_140097944041960: core_fifo_inputs_t;
        signal fifo_full_140097944041960: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944041960: core_fifo_inputs_t;
        signal outputs_full_140097944041960: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944041904: core_fifo_inputs_t;
        signal fifo_full_140097944041904: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944041904: core_fifo_inputs_t;
        signal outputs_full_140097944041904: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944042128: core_fifo_inputs_t;
        signal fifo_full_140097944042128: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944042128: core_fifo_inputs_t;
        signal outputs_full_140097944042128: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944042072: core_fifo_inputs_t;
        signal fifo_full_140097944042072: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944042072: core_fifo_inputs_t;
        signal outputs_full_140097944042072: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944042184: core_fifo_inputs_t;
        signal fifo_full_140097944042184: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944042184: core_fifo_inputs_t;
        signal outputs_full_140097944042184: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944042240: core_fifo_inputs_t;
        signal fifo_full_140097944042240: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944042240: core_fifo_inputs_t;
        signal outputs_full_140097944042240: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944042296: core_fifo_inputs_t;
        signal fifo_full_140097944042296: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944042296: core_fifo_inputs_t;
        signal outputs_full_140097944042296: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944042352: core_fifo_inputs_t;
        signal fifo_full_140097944042352: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944042352: core_fifo_inputs_t;
        signal outputs_full_140097944042352: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944042408: core_fifo_inputs_t;
        signal fifo_full_140097944042408: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944042408: core_fifo_inputs_t;
        signal outputs_full_140097944042408: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944042464: core_fifo_inputs_t;
        signal fifo_full_140097944042464: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944042464: core_fifo_inputs_t;
        signal outputs_full_140097944042464: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944042016: core_fifo_inputs_t;
        signal fifo_full_140097944042016: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944042016: core_fifo_inputs_t;
        signal outputs_full_140097944042016: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944042520: core_fifo_inputs_t;
        signal fifo_full_140097944042520: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944042520: core_fifo_inputs_t;
        signal outputs_full_140097944042520: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944042576: core_fifo_inputs_t;
        signal fifo_full_140097944042576: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944042576: core_fifo_inputs_t;
        signal outputs_full_140097944042576: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944042632: core_fifo_inputs_t;
        signal fifo_full_140097944042632: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944042632: core_fifo_inputs_t;
        signal outputs_full_140097944042632: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944042688: core_fifo_inputs_t;
        signal fifo_full_140097944042688: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944042688: core_fifo_inputs_t;
        signal outputs_full_140097944042688: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944042744: core_fifo_inputs_t;
        signal fifo_full_140097944042744: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944042744: core_fifo_inputs_t;
        signal outputs_full_140097944042744: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944042800: core_fifo_inputs_t;
        signal fifo_full_140097944042800: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944042800: core_fifo_inputs_t;
        signal outputs_full_140097944042800: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944042856: core_fifo_inputs_t;
        signal fifo_full_140097944042856: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944042856: core_fifo_inputs_t;
        signal outputs_full_140097944042856: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944042912: core_fifo_inputs_t;
        signal fifo_full_140097944042912: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944042912: core_fifo_inputs_t;
        signal outputs_full_140097944042912: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944042968: core_fifo_inputs_t;
        signal fifo_full_140097944042968: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944042968: core_fifo_inputs_t;
        signal outputs_full_140097944042968: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944043024: core_fifo_inputs_t;
        signal fifo_full_140097944043024: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944043024: core_fifo_inputs_t;
        signal outputs_full_140097944043024: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944043080: core_fifo_inputs_t;
        signal fifo_full_140097944043080: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944043080: core_fifo_inputs_t;
        signal outputs_full_140097944043080: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944043136: core_fifo_inputs_t;
        signal fifo_full_140097944043136: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944043136: core_fifo_inputs_t;
        signal outputs_full_140097944043136: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944043192: core_fifo_inputs_t;
        signal fifo_full_140097944043192: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944043192: core_fifo_inputs_t;
        signal outputs_full_140097944043192: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944043248: core_fifo_inputs_t;
        signal fifo_full_140097944043248: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944043248: core_fifo_inputs_t;
        signal outputs_full_140097944043248: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944043304: core_fifo_inputs_t;
        signal fifo_full_140097944043304: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944043304: core_fifo_inputs_t;
        signal outputs_full_140097944043304: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944043360: core_fifo_inputs_t;
        signal fifo_full_140097944043360: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944043360: core_fifo_inputs_t;
        signal outputs_full_140097944043360: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944043416: core_fifo_inputs_t;
        signal fifo_full_140097944043416: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944043416: core_fifo_inputs_t;
        signal outputs_full_140097944043416: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944043472: core_fifo_inputs_t;
        signal fifo_full_140097944043472: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944043472: core_fifo_inputs_t;
        signal outputs_full_140097944043472: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944076360: core_fifo_inputs_t;
        signal fifo_full_140097944076360: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944076360: core_fifo_inputs_t;
        signal outputs_full_140097944076360: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944076416: core_fifo_inputs_t;
        signal fifo_full_140097944076416: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944076416: core_fifo_inputs_t;
        signal outputs_full_140097944076416: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944076472: core_fifo_inputs_t;
        signal fifo_full_140097944076472: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944076472: core_fifo_inputs_t;
        signal outputs_full_140097944076472: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944076528: core_fifo_inputs_t;
        signal fifo_full_140097944076528: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944076528: core_fifo_inputs_t;
        signal outputs_full_140097944076528: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944076584: core_fifo_inputs_t;
        signal fifo_full_140097944076584: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944076584: core_fifo_inputs_t;
        signal outputs_full_140097944076584: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944076640: core_fifo_inputs_t;
        signal fifo_full_140097944076640: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944076640: core_fifo_inputs_t;
        signal outputs_full_140097944076640: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944076696: core_fifo_inputs_t;
        signal fifo_full_140097944076696: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944076696: core_fifo_inputs_t;
        signal outputs_full_140097944076696: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944076752: core_fifo_inputs_t;
        signal fifo_full_140097944076752: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944076752: core_fifo_inputs_t;
        signal outputs_full_140097944076752: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944076808: core_fifo_inputs_t;
        signal fifo_full_140097944076808: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944076808: core_fifo_inputs_t;
        signal outputs_full_140097944076808: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944076864: core_fifo_inputs_t;
        signal fifo_full_140097944076864: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944076864: core_fifo_inputs_t;
        signal outputs_full_140097944076864: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944076920: core_fifo_inputs_t;
        signal fifo_full_140097944076920: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944076920: core_fifo_inputs_t;
        signal outputs_full_140097944076920: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944076976: core_fifo_inputs_t;
        signal fifo_full_140097944076976: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944076976: core_fifo_inputs_t;
        signal outputs_full_140097944076976: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944077032: core_fifo_inputs_t;
        signal fifo_full_140097944077032: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944077032: core_fifo_inputs_t;
        signal outputs_full_140097944077032: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944077088: core_fifo_inputs_t;
        signal fifo_full_140097944077088: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944077088: core_fifo_inputs_t;
        signal outputs_full_140097944077088: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944077144: core_fifo_inputs_t;
        signal fifo_full_140097944077144: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944077144: core_fifo_inputs_t;
        signal outputs_full_140097944077144: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944077200: core_fifo_inputs_t;
        signal fifo_full_140097944077200: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944077200: core_fifo_inputs_t;
        signal outputs_full_140097944077200: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944077256: core_fifo_inputs_t;
        signal fifo_full_140097944077256: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944077256: core_fifo_inputs_t;
        signal outputs_full_140097944077256: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944077312: core_fifo_inputs_t;
        signal fifo_full_140097944077312: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944077312: core_fifo_inputs_t;
        signal outputs_full_140097944077312: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944077368: core_fifo_inputs_t;
        signal fifo_full_140097944077368: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944077368: core_fifo_inputs_t;
        signal outputs_full_140097944077368: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944077424: core_fifo_inputs_t;
        signal fifo_full_140097944077424: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944077424: core_fifo_inputs_t;
        signal outputs_full_140097944077424: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944077480: core_fifo_inputs_t;
        signal fifo_full_140097944077480: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944077480: core_fifo_inputs_t;
        signal outputs_full_140097944077480: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944077536: core_fifo_inputs_t;
        signal fifo_full_140097944077536: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944077536: core_fifo_inputs_t;
        signal outputs_full_140097944077536: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944077592: core_fifo_inputs_t;
        signal fifo_full_140097944077592: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944077592: core_fifo_inputs_t;
        signal outputs_full_140097944077592: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944077648: core_fifo_inputs_t;
        signal fifo_full_140097944077648: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944077648: core_fifo_inputs_t;
        signal outputs_full_140097944077648: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944077704: core_fifo_inputs_t;
        signal fifo_full_140097944077704: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944077704: core_fifo_inputs_t;
        signal outputs_full_140097944077704: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944077760: core_fifo_inputs_t;
        signal fifo_full_140097944077760: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944077760: core_fifo_inputs_t;
        signal outputs_full_140097944077760: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944077816: core_fifo_inputs_t;
        signal fifo_full_140097944077816: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944077816: core_fifo_inputs_t;
        signal outputs_full_140097944077816: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944077872: core_fifo_inputs_t;
        signal fifo_full_140097944077872: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944077872: core_fifo_inputs_t;
        signal outputs_full_140097944077872: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944077928: core_fifo_inputs_t;
        signal fifo_full_140097944077928: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944077928: core_fifo_inputs_t;
        signal outputs_full_140097944077928: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944077984: core_fifo_inputs_t;
        signal fifo_full_140097944077984: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944077984: core_fifo_inputs_t;
        signal outputs_full_140097944077984: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944078040: core_fifo_inputs_t;
        signal fifo_full_140097944078040: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944078040: core_fifo_inputs_t;
        signal outputs_full_140097944078040: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944078096: core_fifo_inputs_t;
        signal fifo_full_140097944078096: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944078096: core_fifo_inputs_t;
        signal outputs_full_140097944078096: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944078152: core_fifo_inputs_t;
        signal fifo_full_140097944078152: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944078152: core_fifo_inputs_t;
        signal outputs_full_140097944078152: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944078208: core_fifo_inputs_t;
        signal fifo_full_140097944078208: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944078208: core_fifo_inputs_t;
        signal outputs_full_140097944078208: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944078264: core_fifo_inputs_t;
        signal fifo_full_140097944078264: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944078264: core_fifo_inputs_t;
        signal outputs_full_140097944078264: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944078320: core_fifo_inputs_t;
        signal fifo_full_140097944078320: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944078320: core_fifo_inputs_t;
        signal outputs_full_140097944078320: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944078376: core_fifo_inputs_t;
        signal fifo_full_140097944078376: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944078376: core_fifo_inputs_t;
        signal outputs_full_140097944078376: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944078432: core_fifo_inputs_t;
        signal fifo_full_140097944078432: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944078432: core_fifo_inputs_t;
        signal outputs_full_140097944078432: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944078488: core_fifo_inputs_t;
        signal fifo_full_140097944078488: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944078488: core_fifo_inputs_t;
        signal outputs_full_140097944078488: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944078544: core_fifo_inputs_t;
        signal fifo_full_140097944078544: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944078544: core_fifo_inputs_t;
        signal outputs_full_140097944078544: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944078600: core_fifo_inputs_t;
        signal fifo_full_140097944078600: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944078600: core_fifo_inputs_t;
        signal outputs_full_140097944078600: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944078656: core_fifo_inputs_t;
        signal fifo_full_140097944078656: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944078656: core_fifo_inputs_t;
        signal outputs_full_140097944078656: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944078712: core_fifo_inputs_t;
        signal fifo_full_140097944078712: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944078712: core_fifo_inputs_t;
        signal outputs_full_140097944078712: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944078768: core_fifo_inputs_t;
        signal fifo_full_140097944078768: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944078768: core_fifo_inputs_t;
        signal outputs_full_140097944078768: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944078824: core_fifo_inputs_t;
        signal fifo_full_140097944078824: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944078824: core_fifo_inputs_t;
        signal outputs_full_140097944078824: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944078880: core_fifo_inputs_t;
        signal fifo_full_140097944078880: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944078880: core_fifo_inputs_t;
        signal outputs_full_140097944078880: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944078936: core_fifo_inputs_t;
        signal fifo_full_140097944078936: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944078936: core_fifo_inputs_t;
        signal outputs_full_140097944078936: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944078992: core_fifo_inputs_t;
        signal fifo_full_140097944078992: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944078992: core_fifo_inputs_t;
        signal outputs_full_140097944078992: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944079048: core_fifo_inputs_t;
        signal fifo_full_140097944079048: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944079048: core_fifo_inputs_t;
        signal outputs_full_140097944079048: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944079104: core_fifo_inputs_t;
        signal fifo_full_140097944079104: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944079104: core_fifo_inputs_t;
        signal outputs_full_140097944079104: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944079160: core_fifo_inputs_t;
        signal fifo_full_140097944079160: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944079160: core_fifo_inputs_t;
        signal outputs_full_140097944079160: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944079216: core_fifo_inputs_t;
        signal fifo_full_140097944079216: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944079216: core_fifo_inputs_t;
        signal outputs_full_140097944079216: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944079272: core_fifo_inputs_t;
        signal fifo_full_140097944079272: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944079272: core_fifo_inputs_t;
        signal outputs_full_140097944079272: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944079328: core_fifo_inputs_t;
        signal fifo_full_140097944079328: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944079328: core_fifo_inputs_t;
        signal outputs_full_140097944079328: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944079384: core_fifo_inputs_t;
        signal fifo_full_140097944079384: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944079384: core_fifo_inputs_t;
        signal outputs_full_140097944079384: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944079440: core_fifo_inputs_t;
        signal fifo_full_140097944079440: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944079440: core_fifo_inputs_t;
        signal outputs_full_140097944079440: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944079496: core_fifo_inputs_t;
        signal fifo_full_140097944079496: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944079496: core_fifo_inputs_t;
        signal outputs_full_140097944079496: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944079552: core_fifo_inputs_t;
        signal fifo_full_140097944079552: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944079552: core_fifo_inputs_t;
        signal outputs_full_140097944079552: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944079608: core_fifo_inputs_t;
        signal fifo_full_140097944079608: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944079608: core_fifo_inputs_t;
        signal outputs_full_140097944079608: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944079664: core_fifo_inputs_t;
        signal fifo_full_140097944079664: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944079664: core_fifo_inputs_t;
        signal outputs_full_140097944079664: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944079720: core_fifo_inputs_t;
        signal fifo_full_140097944079720: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944079720: core_fifo_inputs_t;
        signal outputs_full_140097944079720: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944079776: core_fifo_inputs_t;
        signal fifo_full_140097944079776: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944079776: core_fifo_inputs_t;
        signal outputs_full_140097944079776: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944079832: core_fifo_inputs_t;
        signal fifo_full_140097944079832: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944079832: core_fifo_inputs_t;
        signal outputs_full_140097944079832: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944079888: core_fifo_inputs_t;
        signal fifo_full_140097944079888: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944079888: core_fifo_inputs_t;
        signal outputs_full_140097944079888: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944079944: core_fifo_inputs_t;
        signal fifo_full_140097944079944: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944079944: core_fifo_inputs_t;
        signal outputs_full_140097944079944: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944080000: core_fifo_inputs_t;
        signal fifo_full_140097944080000: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944080000: core_fifo_inputs_t;
        signal outputs_full_140097944080000: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944080056: core_fifo_inputs_t;
        signal fifo_full_140097944080056: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944080056: core_fifo_inputs_t;
        signal outputs_full_140097944080056: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944080112: core_fifo_inputs_t;
        signal fifo_full_140097944080112: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944080112: core_fifo_inputs_t;
        signal outputs_full_140097944080112: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944080168: core_fifo_inputs_t;
        signal fifo_full_140097944080168: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944080168: core_fifo_inputs_t;
        signal outputs_full_140097944080168: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944080224: core_fifo_inputs_t;
        signal fifo_full_140097944080224: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944080224: core_fifo_inputs_t;
        signal outputs_full_140097944080224: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944080280: core_fifo_inputs_t;
        signal fifo_full_140097944080280: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944080280: core_fifo_inputs_t;
        signal outputs_full_140097944080280: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944080336: core_fifo_inputs_t;
        signal fifo_full_140097944080336: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944080336: core_fifo_inputs_t;
        signal outputs_full_140097944080336: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944096840: core_fifo_inputs_t;
        signal fifo_full_140097944096840: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944096840: core_fifo_inputs_t;
        signal outputs_full_140097944096840: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944096896: core_fifo_inputs_t;
        signal fifo_full_140097944096896: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944096896: core_fifo_inputs_t;
        signal outputs_full_140097944096896: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944096952: core_fifo_inputs_t;
        signal fifo_full_140097944096952: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944096952: core_fifo_inputs_t;
        signal outputs_full_140097944096952: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944097008: core_fifo_inputs_t;
        signal fifo_full_140097944097008: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944097008: core_fifo_inputs_t;
        signal outputs_full_140097944097008: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944097064: core_fifo_inputs_t;
        signal fifo_full_140097944097064: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944097064: core_fifo_inputs_t;
        signal outputs_full_140097944097064: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944097120: core_fifo_inputs_t;
        signal fifo_full_140097944097120: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944097120: core_fifo_inputs_t;
        signal outputs_full_140097944097120: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944097176: core_fifo_inputs_t;
        signal fifo_full_140097944097176: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944097176: core_fifo_inputs_t;
        signal outputs_full_140097944097176: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944097232: core_fifo_inputs_t;
        signal fifo_full_140097944097232: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944097232: core_fifo_inputs_t;
        signal outputs_full_140097944097232: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944097288: core_fifo_inputs_t;
        signal fifo_full_140097944097288: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944097288: core_fifo_inputs_t;
        signal outputs_full_140097944097288: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944097344: core_fifo_inputs_t;
        signal fifo_full_140097944097344: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944097344: core_fifo_inputs_t;
        signal outputs_full_140097944097344: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944097400: core_fifo_inputs_t;
        signal fifo_full_140097944097400: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944097400: core_fifo_inputs_t;
        signal outputs_full_140097944097400: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944097456: core_fifo_inputs_t;
        signal fifo_full_140097944097456: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944097456: core_fifo_inputs_t;
        signal outputs_full_140097944097456: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944097512: core_fifo_inputs_t;
        signal fifo_full_140097944097512: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944097512: core_fifo_inputs_t;
        signal outputs_full_140097944097512: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944097568: core_fifo_inputs_t;
        signal fifo_full_140097944097568: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944097568: core_fifo_inputs_t;
        signal outputs_full_140097944097568: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944097624: core_fifo_inputs_t;
        signal fifo_full_140097944097624: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944097624: core_fifo_inputs_t;
        signal outputs_full_140097944097624: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944097680: core_fifo_inputs_t;
        signal fifo_full_140097944097680: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944097680: core_fifo_inputs_t;
        signal outputs_full_140097944097680: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944097736: core_fifo_inputs_t;
        signal fifo_full_140097944097736: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944097736: core_fifo_inputs_t;
        signal outputs_full_140097944097736: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944097792: core_fifo_inputs_t;
        signal fifo_full_140097944097792: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944097792: core_fifo_inputs_t;
        signal outputs_full_140097944097792: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944097848: core_fifo_inputs_t;
        signal fifo_full_140097944097848: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944097848: core_fifo_inputs_t;
        signal outputs_full_140097944097848: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944097904: core_fifo_inputs_t;
        signal fifo_full_140097944097904: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944097904: core_fifo_inputs_t;
        signal outputs_full_140097944097904: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944097960: core_fifo_inputs_t;
        signal fifo_full_140097944097960: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944097960: core_fifo_inputs_t;
        signal outputs_full_140097944097960: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944098016: core_fifo_inputs_t;
        signal fifo_full_140097944098016: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944098016: core_fifo_inputs_t;
        signal outputs_full_140097944098016: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944098072: core_fifo_inputs_t;
        signal fifo_full_140097944098072: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944098072: core_fifo_inputs_t;
        signal outputs_full_140097944098072: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944098128: core_fifo_inputs_t;
        signal fifo_full_140097944098128: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944098128: core_fifo_inputs_t;
        signal outputs_full_140097944098128: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944098184: core_fifo_inputs_t;
        signal fifo_full_140097944098184: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944098184: core_fifo_inputs_t;
        signal outputs_full_140097944098184: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944098240: core_fifo_inputs_t;
        signal fifo_full_140097944098240: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944098240: core_fifo_inputs_t;
        signal outputs_full_140097944098240: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944098296: core_fifo_inputs_t;
        signal fifo_full_140097944098296: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944098296: core_fifo_inputs_t;
        signal outputs_full_140097944098296: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944098352: core_fifo_inputs_t;
        signal fifo_full_140097944098352: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944098352: core_fifo_inputs_t;
        signal outputs_full_140097944098352: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944098408: core_fifo_inputs_t;
        signal fifo_full_140097944098408: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944098408: core_fifo_inputs_t;
        signal outputs_full_140097944098408: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944098464: core_fifo_inputs_t;
        signal fifo_full_140097944098464: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944098464: core_fifo_inputs_t;
        signal outputs_full_140097944098464: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944098520: core_fifo_inputs_t;
        signal fifo_full_140097944098520: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944098520: core_fifo_inputs_t;
        signal outputs_full_140097944098520: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944098576: core_fifo_inputs_t;
        signal fifo_full_140097944098576: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944098576: core_fifo_inputs_t;
        signal outputs_full_140097944098576: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944098632: core_fifo_inputs_t;
        signal fifo_full_140097944098632: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944098632: core_fifo_inputs_t;
        signal outputs_full_140097944098632: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944098688: core_fifo_inputs_t;
        signal fifo_full_140097944098688: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944098688: core_fifo_inputs_t;
        signal outputs_full_140097944098688: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944098744: core_fifo_inputs_t;
        signal fifo_full_140097944098744: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944098744: core_fifo_inputs_t;
        signal outputs_full_140097944098744: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944098800: core_fifo_inputs_t;
        signal fifo_full_140097944098800: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944098800: core_fifo_inputs_t;
        signal outputs_full_140097944098800: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944098856: core_fifo_inputs_t;
        signal fifo_full_140097944098856: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944098856: core_fifo_inputs_t;
        signal outputs_full_140097944098856: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944098912: core_fifo_inputs_t;
        signal fifo_full_140097944098912: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944098912: core_fifo_inputs_t;
        signal outputs_full_140097944098912: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944098968: core_fifo_inputs_t;
        signal fifo_full_140097944098968: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944098968: core_fifo_inputs_t;
        signal outputs_full_140097944098968: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944099024: core_fifo_inputs_t;
        signal fifo_full_140097944099024: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944099024: core_fifo_inputs_t;
        signal outputs_full_140097944099024: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944099080: core_fifo_inputs_t;
        signal fifo_full_140097944099080: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944099080: core_fifo_inputs_t;
        signal outputs_full_140097944099080: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944099136: core_fifo_inputs_t;
        signal fifo_full_140097944099136: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944099136: core_fifo_inputs_t;
        signal outputs_full_140097944099136: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944099192: core_fifo_inputs_t;
        signal fifo_full_140097944099192: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944099192: core_fifo_inputs_t;
        signal outputs_full_140097944099192: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944099248: core_fifo_inputs_t;
        signal fifo_full_140097944099248: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944099248: core_fifo_inputs_t;
        signal outputs_full_140097944099248: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944099304: core_fifo_inputs_t;
        signal fifo_full_140097944099304: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944099304: core_fifo_inputs_t;
        signal outputs_full_140097944099304: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944099360: core_fifo_inputs_t;
        signal fifo_full_140097944099360: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944099360: core_fifo_inputs_t;
        signal outputs_full_140097944099360: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944099416: core_fifo_inputs_t;
        signal fifo_full_140097944099416: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944099416: core_fifo_inputs_t;
        signal outputs_full_140097944099416: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944099472: core_fifo_inputs_t;
        signal fifo_full_140097944099472: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944099472: core_fifo_inputs_t;
        signal outputs_full_140097944099472: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944099528: core_fifo_inputs_t;
        signal fifo_full_140097944099528: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944099528: core_fifo_inputs_t;
        signal outputs_full_140097944099528: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097965543496: core_fifo_inputs_t;
        signal fifo_full_140097965543496: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097965543496: core_fifo_inputs_t;
        signal outputs_full_140097965543496: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944041736: core_fifo_inputs_t;
        signal fifo_full_140097944041736: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944041736: core_fifo_inputs_t;
        signal outputs_full_140097944041736: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944041624: core_fifo_inputs_t;
        signal fifo_full_140097944041624: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944041624: core_fifo_inputs_t;
        signal outputs_full_140097944041624: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944041568: core_fifo_inputs_t;
        signal fifo_full_140097944041568: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944041568: core_fifo_inputs_t;
        signal outputs_full_140097944041568: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944041792: core_fifo_inputs_t;
        signal fifo_full_140097944041792: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944041792: core_fifo_inputs_t;
        signal outputs_full_140097944041792: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944041456: core_fifo_inputs_t;
        signal fifo_full_140097944041456: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944041456: core_fifo_inputs_t;
        signal outputs_full_140097944041456: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944099584: core_fifo_inputs_t;
        signal fifo_full_140097944099584: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944099584: core_fifo_inputs_t;
        signal outputs_full_140097944099584: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944099640: core_fifo_inputs_t;
        signal fifo_full_140097944099640: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944099640: core_fifo_inputs_t;
        signal outputs_full_140097944099640: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944099696: core_fifo_inputs_t;
        signal fifo_full_140097944099696: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944099696: core_fifo_inputs_t;
        signal outputs_full_140097944099696: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944099752: core_fifo_inputs_t;
        signal fifo_full_140097944099752: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944099752: core_fifo_inputs_t;
        signal outputs_full_140097944099752: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944099808: core_fifo_inputs_t;
        signal fifo_full_140097944099808: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944099808: core_fifo_inputs_t;
        signal outputs_full_140097944099808: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944099864: core_fifo_inputs_t;
        signal fifo_full_140097944099864: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944099864: core_fifo_inputs_t;
        signal outputs_full_140097944099864: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944099920: core_fifo_inputs_t;
        signal fifo_full_140097944099920: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944099920: core_fifo_inputs_t;
        signal outputs_full_140097944099920: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944099976: core_fifo_inputs_t;
        signal fifo_full_140097944099976: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944099976: core_fifo_inputs_t;
        signal outputs_full_140097944099976: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944100032: core_fifo_inputs_t;
        signal fifo_full_140097944100032: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944100032: core_fifo_inputs_t;
        signal outputs_full_140097944100032: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944100088: core_fifo_inputs_t;
        signal fifo_full_140097944100088: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944100088: core_fifo_inputs_t;
        signal outputs_full_140097944100088: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944100144: core_fifo_inputs_t;
        signal fifo_full_140097944100144: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944100144: core_fifo_inputs_t;
        signal outputs_full_140097944100144: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944100200: core_fifo_inputs_t;
        signal fifo_full_140097944100200: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944100200: core_fifo_inputs_t;
        signal outputs_full_140097944100200: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944100256: core_fifo_inputs_t;
        signal fifo_full_140097944100256: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944100256: core_fifo_inputs_t;
        signal outputs_full_140097944100256: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944100312: core_fifo_inputs_t;
        signal fifo_full_140097944100312: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944100312: core_fifo_inputs_t;
        signal outputs_full_140097944100312: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944100368: core_fifo_inputs_t;
        signal fifo_full_140097944100368: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944100368: core_fifo_inputs_t;
        signal outputs_full_140097944100368: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944100424: core_fifo_inputs_t;
        signal fifo_full_140097944100424: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944100424: core_fifo_inputs_t;
        signal outputs_full_140097944100424: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944100480: core_fifo_inputs_t;
        signal fifo_full_140097944100480: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944100480: core_fifo_inputs_t;
        signal outputs_full_140097944100480: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944100536: core_fifo_inputs_t;
        signal fifo_full_140097944100536: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944100536: core_fifo_inputs_t;
        signal outputs_full_140097944100536: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944100592: core_fifo_inputs_t;
        signal fifo_full_140097944100592: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944100592: core_fifo_inputs_t;
        signal outputs_full_140097944100592: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944100648: core_fifo_inputs_t;
        signal fifo_full_140097944100648: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944100648: core_fifo_inputs_t;
        signal outputs_full_140097944100648: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944100704: core_fifo_inputs_t;
        signal fifo_full_140097944100704: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944100704: core_fifo_inputs_t;
        signal outputs_full_140097944100704: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944100760: core_fifo_inputs_t;
        signal fifo_full_140097944100760: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944100760: core_fifo_inputs_t;
        signal outputs_full_140097944100760: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944100816: core_fifo_inputs_t;
        signal fifo_full_140097944100816: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944100816: core_fifo_inputs_t;
        signal outputs_full_140097944100816: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944113224: core_fifo_inputs_t;
        signal fifo_full_140097944113224: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944113224: core_fifo_inputs_t;
        signal outputs_full_140097944113224: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944113280: core_fifo_inputs_t;
        signal fifo_full_140097944113280: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944113280: core_fifo_inputs_t;
        signal outputs_full_140097944113280: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944113336: core_fifo_inputs_t;
        signal fifo_full_140097944113336: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944113336: core_fifo_inputs_t;
        signal outputs_full_140097944113336: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944113392: core_fifo_inputs_t;
        signal fifo_full_140097944113392: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944113392: core_fifo_inputs_t;
        signal outputs_full_140097944113392: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944113448: core_fifo_inputs_t;
        signal fifo_full_140097944113448: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944113448: core_fifo_inputs_t;
        signal outputs_full_140097944113448: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944113504: core_fifo_inputs_t;
        signal fifo_full_140097944113504: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944113504: core_fifo_inputs_t;
        signal outputs_full_140097944113504: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944113560: core_fifo_inputs_t;
        signal fifo_full_140097944113560: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944113560: core_fifo_inputs_t;
        signal outputs_full_140097944113560: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944113616: core_fifo_inputs_t;
        signal fifo_full_140097944113616: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944113616: core_fifo_inputs_t;
        signal outputs_full_140097944113616: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944113672: core_fifo_inputs_t;
        signal fifo_full_140097944113672: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944113672: core_fifo_inputs_t;
        signal outputs_full_140097944113672: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944113728: core_fifo_inputs_t;
        signal fifo_full_140097944113728: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944113728: core_fifo_inputs_t;
        signal outputs_full_140097944113728: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944113784: core_fifo_inputs_t;
        signal fifo_full_140097944113784: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944113784: core_fifo_inputs_t;
        signal outputs_full_140097944113784: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944113840: core_fifo_inputs_t;
        signal fifo_full_140097944113840: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944113840: core_fifo_inputs_t;
        signal outputs_full_140097944113840: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944113896: core_fifo_inputs_t;
        signal fifo_full_140097944113896: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944113896: core_fifo_inputs_t;
        signal outputs_full_140097944113896: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944113952: core_fifo_inputs_t;
        signal fifo_full_140097944113952: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944113952: core_fifo_inputs_t;
        signal outputs_full_140097944113952: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944114008: core_fifo_inputs_t;
        signal fifo_full_140097944114008: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944114008: core_fifo_inputs_t;
        signal outputs_full_140097944114008: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944114064: core_fifo_inputs_t;
        signal fifo_full_140097944114064: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944114064: core_fifo_inputs_t;
        signal outputs_full_140097944114064: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944114120: core_fifo_inputs_t;
        signal fifo_full_140097944114120: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944114120: core_fifo_inputs_t;
        signal outputs_full_140097944114120: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944114176: core_fifo_inputs_t;
        signal fifo_full_140097944114176: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944114176: core_fifo_inputs_t;
        signal outputs_full_140097944114176: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944114232: core_fifo_inputs_t;
        signal fifo_full_140097944114232: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944114232: core_fifo_inputs_t;
        signal outputs_full_140097944114232: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944114288: core_fifo_inputs_t;
        signal fifo_full_140097944114288: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944114288: core_fifo_inputs_t;
        signal outputs_full_140097944114288: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944114344: core_fifo_inputs_t;
        signal fifo_full_140097944114344: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944114344: core_fifo_inputs_t;
        signal outputs_full_140097944114344: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944114400: core_fifo_inputs_t;
        signal fifo_full_140097944114400: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944114400: core_fifo_inputs_t;
        signal outputs_full_140097944114400: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944114456: core_fifo_inputs_t;
        signal fifo_full_140097944114456: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944114456: core_fifo_inputs_t;
        signal outputs_full_140097944114456: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944114512: core_fifo_inputs_t;
        signal fifo_full_140097944114512: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944114512: core_fifo_inputs_t;
        signal outputs_full_140097944114512: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944114568: core_fifo_inputs_t;
        signal fifo_full_140097944114568: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944114568: core_fifo_inputs_t;
        signal outputs_full_140097944114568: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944114624: core_fifo_inputs_t;
        signal fifo_full_140097944114624: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944114624: core_fifo_inputs_t;
        signal outputs_full_140097944114624: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944114680: core_fifo_inputs_t;
        signal fifo_full_140097944114680: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944114680: core_fifo_inputs_t;
        signal outputs_full_140097944114680: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944114736: core_fifo_inputs_t;
        signal fifo_full_140097944114736: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944114736: core_fifo_inputs_t;
        signal outputs_full_140097944114736: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944114792: core_fifo_inputs_t;
        signal fifo_full_140097944114792: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944114792: core_fifo_inputs_t;
        signal outputs_full_140097944114792: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944114848: core_fifo_inputs_t;
        signal fifo_full_140097944114848: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944114848: core_fifo_inputs_t;
        signal outputs_full_140097944114848: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944114904: core_fifo_inputs_t;
        signal fifo_full_140097944114904: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944114904: core_fifo_inputs_t;
        signal outputs_full_140097944114904: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944114960: core_fifo_inputs_t;
        signal fifo_full_140097944114960: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944114960: core_fifo_inputs_t;
        signal outputs_full_140097944114960: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944115016: core_fifo_inputs_t;
        signal fifo_full_140097944115016: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944115016: core_fifo_inputs_t;
        signal outputs_full_140097944115016: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944115072: core_fifo_inputs_t;
        signal fifo_full_140097944115072: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944115072: core_fifo_inputs_t;
        signal outputs_full_140097944115072: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944115128: core_fifo_inputs_t;
        signal fifo_full_140097944115128: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944115128: core_fifo_inputs_t;
        signal outputs_full_140097944115128: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944115184: core_fifo_inputs_t;
        signal fifo_full_140097944115184: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944115184: core_fifo_inputs_t;
        signal outputs_full_140097944115184: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944115240: core_fifo_inputs_t;
        signal fifo_full_140097944115240: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944115240: core_fifo_inputs_t;
        signal outputs_full_140097944115240: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944115296: core_fifo_inputs_t;
        signal fifo_full_140097944115296: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944115296: core_fifo_inputs_t;
        signal outputs_full_140097944115296: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944115352: core_fifo_inputs_t;
        signal fifo_full_140097944115352: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944115352: core_fifo_inputs_t;
        signal outputs_full_140097944115352: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944115408: core_fifo_inputs_t;
        signal fifo_full_140097944115408: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944115408: core_fifo_inputs_t;
        signal outputs_full_140097944115408: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944115464: core_fifo_inputs_t;
        signal fifo_full_140097944115464: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944115464: core_fifo_inputs_t;
        signal outputs_full_140097944115464: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944115520: core_fifo_inputs_t;
        signal fifo_full_140097944115520: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944115520: core_fifo_inputs_t;
        signal outputs_full_140097944115520: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944115576: core_fifo_inputs_t;
        signal fifo_full_140097944115576: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944115576: core_fifo_inputs_t;
        signal outputs_full_140097944115576: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944115632: core_fifo_inputs_t;
        signal fifo_full_140097944115632: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944115632: core_fifo_inputs_t;
        signal outputs_full_140097944115632: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944115688: core_fifo_inputs_t;
        signal fifo_full_140097944115688: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944115688: core_fifo_inputs_t;
        signal outputs_full_140097944115688: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944115744: core_fifo_inputs_t;
        signal fifo_full_140097944115744: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944115744: core_fifo_inputs_t;
        signal outputs_full_140097944115744: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944115800: core_fifo_inputs_t;
        signal fifo_full_140097944115800: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944115800: core_fifo_inputs_t;
        signal outputs_full_140097944115800: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944115856: core_fifo_inputs_t;
        signal fifo_full_140097944115856: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944115856: core_fifo_inputs_t;
        signal outputs_full_140097944115856: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944115912: core_fifo_inputs_t;
        signal fifo_full_140097944115912: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944115912: core_fifo_inputs_t;
        signal outputs_full_140097944115912: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944115968: core_fifo_inputs_t;
        signal fifo_full_140097944115968: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944115968: core_fifo_inputs_t;
        signal outputs_full_140097944115968: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944116024: core_fifo_inputs_t;
        signal fifo_full_140097944116024: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944116024: core_fifo_inputs_t;
        signal outputs_full_140097944116024: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944116080: core_fifo_inputs_t;
        signal fifo_full_140097944116080: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944116080: core_fifo_inputs_t;
        signal outputs_full_140097944116080: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944116136: core_fifo_inputs_t;
        signal fifo_full_140097944116136: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944116136: core_fifo_inputs_t;
        signal outputs_full_140097944116136: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944116192: core_fifo_inputs_t;
        signal fifo_full_140097944116192: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944116192: core_fifo_inputs_t;
        signal outputs_full_140097944116192: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944116248: core_fifo_inputs_t;
        signal fifo_full_140097944116248: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944116248: core_fifo_inputs_t;
        signal outputs_full_140097944116248: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944116304: core_fifo_inputs_t;
        signal fifo_full_140097944116304: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944116304: core_fifo_inputs_t;
        signal outputs_full_140097944116304: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944116360: core_fifo_inputs_t;
        signal fifo_full_140097944116360: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944116360: core_fifo_inputs_t;
        signal outputs_full_140097944116360: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944116416: core_fifo_inputs_t;
        signal fifo_full_140097944116416: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944116416: core_fifo_inputs_t;
        signal outputs_full_140097944116416: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944116472: core_fifo_inputs_t;
        signal fifo_full_140097944116472: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944116472: core_fifo_inputs_t;
        signal outputs_full_140097944116472: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944116528: core_fifo_inputs_t;
        signal fifo_full_140097944116528: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944116528: core_fifo_inputs_t;
        signal outputs_full_140097944116528: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944116584: core_fifo_inputs_t;
        signal fifo_full_140097944116584: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944116584: core_fifo_inputs_t;
        signal outputs_full_140097944116584: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944116640: core_fifo_inputs_t;
        signal fifo_full_140097944116640: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944116640: core_fifo_inputs_t;
        signal outputs_full_140097944116640: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944116696: core_fifo_inputs_t;
        signal fifo_full_140097944116696: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944116696: core_fifo_inputs_t;
        signal outputs_full_140097944116696: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944116752: core_fifo_inputs_t;
        signal fifo_full_140097944116752: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944116752: core_fifo_inputs_t;
        signal outputs_full_140097944116752: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944116808: core_fifo_inputs_t;
        signal fifo_full_140097944116808: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944116808: core_fifo_inputs_t;
        signal outputs_full_140097944116808: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944116864: core_fifo_inputs_t;
        signal fifo_full_140097944116864: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944116864: core_fifo_inputs_t;
        signal outputs_full_140097944116864: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944116920: core_fifo_inputs_t;
        signal fifo_full_140097944116920: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944116920: core_fifo_inputs_t;
        signal outputs_full_140097944116920: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944116976: core_fifo_inputs_t;
        signal fifo_full_140097944116976: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944116976: core_fifo_inputs_t;
        signal outputs_full_140097944116976: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944117032: core_fifo_inputs_t;
        signal fifo_full_140097944117032: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944117032: core_fifo_inputs_t;
        signal outputs_full_140097944117032: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944117088: core_fifo_inputs_t;
        signal fifo_full_140097944117088: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944117088: core_fifo_inputs_t;
        signal outputs_full_140097944117088: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944117144: core_fifo_inputs_t;
        signal fifo_full_140097944117144: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944117144: core_fifo_inputs_t;
        signal outputs_full_140097944117144: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944117200: core_fifo_inputs_t;
        signal fifo_full_140097944117200: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944117200: core_fifo_inputs_t;
        signal outputs_full_140097944117200: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944125512: core_fifo_inputs_t;
        signal fifo_full_140097944125512: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944125512: core_fifo_inputs_t;
        signal outputs_full_140097944125512: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944125568: core_fifo_inputs_t;
        signal fifo_full_140097944125568: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944125568: core_fifo_inputs_t;
        signal outputs_full_140097944125568: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944125624: core_fifo_inputs_t;
        signal fifo_full_140097944125624: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944125624: core_fifo_inputs_t;
        signal outputs_full_140097944125624: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944125680: core_fifo_inputs_t;
        signal fifo_full_140097944125680: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944125680: core_fifo_inputs_t;
        signal outputs_full_140097944125680: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944125736: core_fifo_inputs_t;
        signal fifo_full_140097944125736: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944125736: core_fifo_inputs_t;
        signal outputs_full_140097944125736: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944125792: core_fifo_inputs_t;
        signal fifo_full_140097944125792: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944125792: core_fifo_inputs_t;
        signal outputs_full_140097944125792: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944125848: core_fifo_inputs_t;
        signal fifo_full_140097944125848: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944125848: core_fifo_inputs_t;
        signal outputs_full_140097944125848: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944125904: core_fifo_inputs_t;
        signal fifo_full_140097944125904: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944125904: core_fifo_inputs_t;
        signal outputs_full_140097944125904: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944125960: core_fifo_inputs_t;
        signal fifo_full_140097944125960: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944125960: core_fifo_inputs_t;
        signal outputs_full_140097944125960: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944126016: core_fifo_inputs_t;
        signal fifo_full_140097944126016: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944126016: core_fifo_inputs_t;
        signal outputs_full_140097944126016: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944126072: core_fifo_inputs_t;
        signal fifo_full_140097944126072: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944126072: core_fifo_inputs_t;
        signal outputs_full_140097944126072: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944126128: core_fifo_inputs_t;
        signal fifo_full_140097944126128: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944126128: core_fifo_inputs_t;
        signal outputs_full_140097944126128: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944126184: core_fifo_inputs_t;
        signal fifo_full_140097944126184: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944126184: core_fifo_inputs_t;
        signal outputs_full_140097944126184: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944126240: core_fifo_inputs_t;
        signal fifo_full_140097944126240: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944126240: core_fifo_inputs_t;
        signal outputs_full_140097944126240: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944126296: core_fifo_inputs_t;
        signal fifo_full_140097944126296: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944126296: core_fifo_inputs_t;
        signal outputs_full_140097944126296: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944126352: core_fifo_inputs_t;
        signal fifo_full_140097944126352: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944126352: core_fifo_inputs_t;
        signal outputs_full_140097944126352: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944126408: core_fifo_inputs_t;
        signal fifo_full_140097944126408: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944126408: core_fifo_inputs_t;
        signal outputs_full_140097944126408: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944126464: core_fifo_inputs_t;
        signal fifo_full_140097944126464: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944126464: core_fifo_inputs_t;
        signal outputs_full_140097944126464: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944126520: core_fifo_inputs_t;
        signal fifo_full_140097944126520: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944126520: core_fifo_inputs_t;
        signal outputs_full_140097944126520: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944126576: core_fifo_inputs_t;
        signal fifo_full_140097944126576: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944126576: core_fifo_inputs_t;
        signal outputs_full_140097944126576: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944126632: core_fifo_inputs_t;
        signal fifo_full_140097944126632: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944126632: core_fifo_inputs_t;
        signal outputs_full_140097944126632: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944126688: core_fifo_inputs_t;
        signal fifo_full_140097944126688: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944126688: core_fifo_inputs_t;
        signal outputs_full_140097944126688: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944126744: core_fifo_inputs_t;
        signal fifo_full_140097944126744: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944126744: core_fifo_inputs_t;
        signal outputs_full_140097944126744: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944126800: core_fifo_inputs_t;
        signal fifo_full_140097944126800: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944126800: core_fifo_inputs_t;
        signal outputs_full_140097944126800: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944126856: core_fifo_inputs_t;
        signal fifo_full_140097944126856: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944126856: core_fifo_inputs_t;
        signal outputs_full_140097944126856: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944126912: core_fifo_inputs_t;
        signal fifo_full_140097944126912: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944126912: core_fifo_inputs_t;
        signal outputs_full_140097944126912: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944126968: core_fifo_inputs_t;
        signal fifo_full_140097944126968: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944126968: core_fifo_inputs_t;
        signal outputs_full_140097944126968: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944127024: core_fifo_inputs_t;
        signal fifo_full_140097944127024: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944127024: core_fifo_inputs_t;
        signal outputs_full_140097944127024: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944127080: core_fifo_inputs_t;
        signal fifo_full_140097944127080: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944127080: core_fifo_inputs_t;
        signal outputs_full_140097944127080: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944127136: core_fifo_inputs_t;
        signal fifo_full_140097944127136: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944127136: core_fifo_inputs_t;
        signal outputs_full_140097944127136: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944127192: core_fifo_inputs_t;
        signal fifo_full_140097944127192: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944127192: core_fifo_inputs_t;
        signal outputs_full_140097944127192: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944127248: core_fifo_inputs_t;
        signal fifo_full_140097944127248: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944127248: core_fifo_inputs_t;
        signal outputs_full_140097944127248: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944127304: core_fifo_inputs_t;
        signal fifo_full_140097944127304: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944127304: core_fifo_inputs_t;
        signal outputs_full_140097944127304: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944127360: core_fifo_inputs_t;
        signal fifo_full_140097944127360: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944127360: core_fifo_inputs_t;
        signal outputs_full_140097944127360: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944127416: core_fifo_inputs_t;
        signal fifo_full_140097944127416: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944127416: core_fifo_inputs_t;
        signal outputs_full_140097944127416: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944127472: core_fifo_inputs_t;
        signal fifo_full_140097944127472: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944127472: core_fifo_inputs_t;
        signal outputs_full_140097944127472: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944127528: core_fifo_inputs_t;
        signal fifo_full_140097944127528: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944127528: core_fifo_inputs_t;
        signal outputs_full_140097944127528: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944127584: core_fifo_inputs_t;
        signal fifo_full_140097944127584: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944127584: core_fifo_inputs_t;
        signal outputs_full_140097944127584: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944127640: core_fifo_inputs_t;
        signal fifo_full_140097944127640: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944127640: core_fifo_inputs_t;
        signal outputs_full_140097944127640: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944127696: core_fifo_inputs_t;
        signal fifo_full_140097944127696: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944127696: core_fifo_inputs_t;
        signal outputs_full_140097944127696: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944127752: core_fifo_inputs_t;
        signal fifo_full_140097944127752: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944127752: core_fifo_inputs_t;
        signal outputs_full_140097944127752: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944127808: core_fifo_inputs_t;
        signal fifo_full_140097944127808: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944127808: core_fifo_inputs_t;
        signal outputs_full_140097944127808: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944127864: core_fifo_inputs_t;
        signal fifo_full_140097944127864: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944127864: core_fifo_inputs_t;
        signal outputs_full_140097944127864: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944127920: core_fifo_inputs_t;
        signal fifo_full_140097944127920: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944127920: core_fifo_inputs_t;
        signal outputs_full_140097944127920: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944127976: core_fifo_inputs_t;
        signal fifo_full_140097944127976: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944127976: core_fifo_inputs_t;
        signal outputs_full_140097944127976: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944128032: core_fifo_inputs_t;
        signal fifo_full_140097944128032: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944128032: core_fifo_inputs_t;
        signal outputs_full_140097944128032: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944128088: core_fifo_inputs_t;
        signal fifo_full_140097944128088: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944128088: core_fifo_inputs_t;
        signal outputs_full_140097944128088: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944128144: core_fifo_inputs_t;
        signal fifo_full_140097944128144: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944128144: core_fifo_inputs_t;
        signal outputs_full_140097944128144: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944128200: core_fifo_inputs_t;
        signal fifo_full_140097944128200: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944128200: core_fifo_inputs_t;
        signal outputs_full_140097944128200: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944128256: core_fifo_inputs_t;
        signal fifo_full_140097944128256: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944128256: core_fifo_inputs_t;
        signal outputs_full_140097944128256: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944128312: core_fifo_inputs_t;
        signal fifo_full_140097944128312: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944128312: core_fifo_inputs_t;
        signal outputs_full_140097944128312: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944128368: core_fifo_inputs_t;
        signal fifo_full_140097944128368: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944128368: core_fifo_inputs_t;
        signal outputs_full_140097944128368: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944128424: core_fifo_inputs_t;
        signal fifo_full_140097944128424: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944128424: core_fifo_inputs_t;
        signal outputs_full_140097944128424: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944128480: core_fifo_inputs_t;
        signal fifo_full_140097944128480: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944128480: core_fifo_inputs_t;
        signal outputs_full_140097944128480: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944128536: core_fifo_inputs_t;
        signal fifo_full_140097944128536: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944128536: core_fifo_inputs_t;
        signal outputs_full_140097944128536: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944128592: core_fifo_inputs_t;
        signal fifo_full_140097944128592: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944128592: core_fifo_inputs_t;
        signal outputs_full_140097944128592: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944128648: core_fifo_inputs_t;
        signal fifo_full_140097944128648: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944128648: core_fifo_inputs_t;
        signal outputs_full_140097944128648: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944128704: core_fifo_inputs_t;
        signal fifo_full_140097944128704: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944128704: core_fifo_inputs_t;
        signal outputs_full_140097944128704: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944128760: core_fifo_inputs_t;
        signal fifo_full_140097944128760: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944128760: core_fifo_inputs_t;
        signal outputs_full_140097944128760: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944128816: core_fifo_inputs_t;
        signal fifo_full_140097944128816: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944128816: core_fifo_inputs_t;
        signal outputs_full_140097944128816: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944128872: core_fifo_inputs_t;
        signal fifo_full_140097944128872: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944128872: core_fifo_inputs_t;
        signal outputs_full_140097944128872: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944128928: core_fifo_inputs_t;
        signal fifo_full_140097944128928: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944128928: core_fifo_inputs_t;
        signal outputs_full_140097944128928: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944128984: core_fifo_inputs_t;
        signal fifo_full_140097944128984: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944128984: core_fifo_inputs_t;
        signal outputs_full_140097944128984: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944129040: core_fifo_inputs_t;
        signal fifo_full_140097944129040: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944129040: core_fifo_inputs_t;
        signal outputs_full_140097944129040: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944129096: core_fifo_inputs_t;
        signal fifo_full_140097944129096: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944129096: core_fifo_inputs_t;
        signal outputs_full_140097944129096: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944129152: core_fifo_inputs_t;
        signal fifo_full_140097944129152: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944129152: core_fifo_inputs_t;
        signal outputs_full_140097944129152: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944129208: core_fifo_inputs_t;
        signal fifo_full_140097944129208: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944129208: core_fifo_inputs_t;
        signal outputs_full_140097944129208: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944129264: core_fifo_inputs_t;
        signal fifo_full_140097944129264: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944129264: core_fifo_inputs_t;
        signal outputs_full_140097944129264: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944129320: core_fifo_inputs_t;
        signal fifo_full_140097944129320: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944129320: core_fifo_inputs_t;
        signal outputs_full_140097944129320: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944129376: core_fifo_inputs_t;
        signal fifo_full_140097944129376: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944129376: core_fifo_inputs_t;
        signal outputs_full_140097944129376: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944129432: core_fifo_inputs_t;
        signal fifo_full_140097944129432: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944129432: core_fifo_inputs_t;
        signal outputs_full_140097944129432: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944129488: core_fifo_inputs_t;
        signal fifo_full_140097944129488: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944129488: core_fifo_inputs_t;
        signal outputs_full_140097944129488: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944141896: core_fifo_inputs_t;
        signal fifo_full_140097944141896: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944141896: core_fifo_inputs_t;
        signal outputs_full_140097944141896: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944141952: core_fifo_inputs_t;
        signal fifo_full_140097944141952: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944141952: core_fifo_inputs_t;
        signal outputs_full_140097944141952: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944142008: core_fifo_inputs_t;
        signal fifo_full_140097944142008: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944142008: core_fifo_inputs_t;
        signal outputs_full_140097944142008: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944142064: core_fifo_inputs_t;
        signal fifo_full_140097944142064: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944142064: core_fifo_inputs_t;
        signal outputs_full_140097944142064: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944142120: core_fifo_inputs_t;
        signal fifo_full_140097944142120: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944142120: core_fifo_inputs_t;
        signal outputs_full_140097944142120: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944142176: core_fifo_inputs_t;
        signal fifo_full_140097944142176: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944142176: core_fifo_inputs_t;
        signal outputs_full_140097944142176: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944142232: core_fifo_inputs_t;
        signal fifo_full_140097944142232: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944142232: core_fifo_inputs_t;
        signal outputs_full_140097944142232: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944142288: core_fifo_inputs_t;
        signal fifo_full_140097944142288: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944142288: core_fifo_inputs_t;
        signal outputs_full_140097944142288: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944142344: core_fifo_inputs_t;
        signal fifo_full_140097944142344: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944142344: core_fifo_inputs_t;
        signal outputs_full_140097944142344: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944142400: core_fifo_inputs_t;
        signal fifo_full_140097944142400: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944142400: core_fifo_inputs_t;
        signal outputs_full_140097944142400: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944142456: core_fifo_inputs_t;
        signal fifo_full_140097944142456: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944142456: core_fifo_inputs_t;
        signal outputs_full_140097944142456: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944142512: core_fifo_inputs_t;
        signal fifo_full_140097944142512: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944142512: core_fifo_inputs_t;
        signal outputs_full_140097944142512: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944142568: core_fifo_inputs_t;
        signal fifo_full_140097944142568: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944142568: core_fifo_inputs_t;
        signal outputs_full_140097944142568: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944142624: core_fifo_inputs_t;
        signal fifo_full_140097944142624: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944142624: core_fifo_inputs_t;
        signal outputs_full_140097944142624: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944142680: core_fifo_inputs_t;
        signal fifo_full_140097944142680: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944142680: core_fifo_inputs_t;
        signal outputs_full_140097944142680: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944142736: core_fifo_inputs_t;
        signal fifo_full_140097944142736: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944142736: core_fifo_inputs_t;
        signal outputs_full_140097944142736: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944142792: core_fifo_inputs_t;
        signal fifo_full_140097944142792: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944142792: core_fifo_inputs_t;
        signal outputs_full_140097944142792: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944142848: core_fifo_inputs_t;
        signal fifo_full_140097944142848: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944142848: core_fifo_inputs_t;
        signal outputs_full_140097944142848: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944142904: core_fifo_inputs_t;
        signal fifo_full_140097944142904: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944142904: core_fifo_inputs_t;
        signal outputs_full_140097944142904: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944142960: core_fifo_inputs_t;
        signal fifo_full_140097944142960: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944142960: core_fifo_inputs_t;
        signal outputs_full_140097944142960: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944143016: core_fifo_inputs_t;
        signal fifo_full_140097944143016: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944143016: core_fifo_inputs_t;
        signal outputs_full_140097944143016: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944143072: core_fifo_inputs_t;
        signal fifo_full_140097944143072: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944143072: core_fifo_inputs_t;
        signal outputs_full_140097944143072: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944143128: core_fifo_inputs_t;
        signal fifo_full_140097944143128: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944143128: core_fifo_inputs_t;
        signal outputs_full_140097944143128: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944143184: core_fifo_inputs_t;
        signal fifo_full_140097944143184: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944143184: core_fifo_inputs_t;
        signal outputs_full_140097944143184: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944143240: core_fifo_inputs_t;
        signal fifo_full_140097944143240: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944143240: core_fifo_inputs_t;
        signal outputs_full_140097944143240: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944143296: core_fifo_inputs_t;
        signal fifo_full_140097944143296: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944143296: core_fifo_inputs_t;
        signal outputs_full_140097944143296: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944143352: core_fifo_inputs_t;
        signal fifo_full_140097944143352: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944143352: core_fifo_inputs_t;
        signal outputs_full_140097944143352: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944143408: core_fifo_inputs_t;
        signal fifo_full_140097944143408: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944143408: core_fifo_inputs_t;
        signal outputs_full_140097944143408: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944143464: core_fifo_inputs_t;
        signal fifo_full_140097944143464: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944143464: core_fifo_inputs_t;
        signal outputs_full_140097944143464: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944143520: core_fifo_inputs_t;
        signal fifo_full_140097944143520: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944143520: core_fifo_inputs_t;
        signal outputs_full_140097944143520: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944143576: core_fifo_inputs_t;
        signal fifo_full_140097944143576: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944143576: core_fifo_inputs_t;
        signal outputs_full_140097944143576: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944143632: core_fifo_inputs_t;
        signal fifo_full_140097944143632: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944143632: core_fifo_inputs_t;
        signal outputs_full_140097944143632: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944143688: core_fifo_inputs_t;
        signal fifo_full_140097944143688: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944143688: core_fifo_inputs_t;
        signal outputs_full_140097944143688: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944143744: core_fifo_inputs_t;
        signal fifo_full_140097944143744: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944143744: core_fifo_inputs_t;
        signal outputs_full_140097944143744: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944143800: core_fifo_inputs_t;
        signal fifo_full_140097944143800: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944143800: core_fifo_inputs_t;
        signal outputs_full_140097944143800: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944143856: core_fifo_inputs_t;
        signal fifo_full_140097944143856: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944143856: core_fifo_inputs_t;
        signal outputs_full_140097944143856: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944143912: core_fifo_inputs_t;
        signal fifo_full_140097944143912: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944143912: core_fifo_inputs_t;
        signal outputs_full_140097944143912: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944143968: core_fifo_inputs_t;
        signal fifo_full_140097944143968: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944143968: core_fifo_inputs_t;
        signal outputs_full_140097944143968: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944144024: core_fifo_inputs_t;
        signal fifo_full_140097944144024: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944144024: core_fifo_inputs_t;
        signal outputs_full_140097944144024: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944144080: core_fifo_inputs_t;
        signal fifo_full_140097944144080: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944144080: core_fifo_inputs_t;
        signal outputs_full_140097944144080: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944144136: core_fifo_inputs_t;
        signal fifo_full_140097944144136: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944144136: core_fifo_inputs_t;
        signal outputs_full_140097944144136: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944144192: core_fifo_inputs_t;
        signal fifo_full_140097944144192: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944144192: core_fifo_inputs_t;
        signal outputs_full_140097944144192: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944144248: core_fifo_inputs_t;
        signal fifo_full_140097944144248: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944144248: core_fifo_inputs_t;
        signal outputs_full_140097944144248: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944144304: core_fifo_inputs_t;
        signal fifo_full_140097944144304: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944144304: core_fifo_inputs_t;
        signal outputs_full_140097944144304: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944144360: core_fifo_inputs_t;
        signal fifo_full_140097944144360: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944144360: core_fifo_inputs_t;
        signal outputs_full_140097944144360: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944144416: core_fifo_inputs_t;
        signal fifo_full_140097944144416: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944144416: core_fifo_inputs_t;
        signal outputs_full_140097944144416: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944144472: core_fifo_inputs_t;
        signal fifo_full_140097944144472: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944144472: core_fifo_inputs_t;
        signal outputs_full_140097944144472: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944144528: core_fifo_inputs_t;
        signal fifo_full_140097944144528: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944144528: core_fifo_inputs_t;
        signal outputs_full_140097944144528: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944144584: core_fifo_inputs_t;
        signal fifo_full_140097944144584: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944144584: core_fifo_inputs_t;
        signal outputs_full_140097944144584: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944144640: core_fifo_inputs_t;
        signal fifo_full_140097944144640: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944144640: core_fifo_inputs_t;
        signal outputs_full_140097944144640: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944144696: core_fifo_inputs_t;
        signal fifo_full_140097944144696: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944144696: core_fifo_inputs_t;
        signal outputs_full_140097944144696: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944144752: core_fifo_inputs_t;
        signal fifo_full_140097944144752: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944144752: core_fifo_inputs_t;
        signal outputs_full_140097944144752: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944144808: core_fifo_inputs_t;
        signal fifo_full_140097944144808: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944144808: core_fifo_inputs_t;
        signal outputs_full_140097944144808: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944144864: core_fifo_inputs_t;
        signal fifo_full_140097944144864: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944144864: core_fifo_inputs_t;
        signal outputs_full_140097944144864: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944144920: core_fifo_inputs_t;
        signal fifo_full_140097944144920: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944144920: core_fifo_inputs_t;
        signal outputs_full_140097944144920: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944144976: core_fifo_inputs_t;
        signal fifo_full_140097944144976: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944144976: core_fifo_inputs_t;
        signal outputs_full_140097944144976: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944145032: core_fifo_inputs_t;
        signal fifo_full_140097944145032: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944145032: core_fifo_inputs_t;
        signal outputs_full_140097944145032: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944145088: core_fifo_inputs_t;
        signal fifo_full_140097944145088: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944145088: core_fifo_inputs_t;
        signal outputs_full_140097944145088: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944145144: core_fifo_inputs_t;
        signal fifo_full_140097944145144: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944145144: core_fifo_inputs_t;
        signal outputs_full_140097944145144: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944145200: core_fifo_inputs_t;
        signal fifo_full_140097944145200: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944145200: core_fifo_inputs_t;
        signal outputs_full_140097944145200: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944145256: core_fifo_inputs_t;
        signal fifo_full_140097944145256: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944145256: core_fifo_inputs_t;
        signal outputs_full_140097944145256: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944145312: core_fifo_inputs_t;
        signal fifo_full_140097944145312: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944145312: core_fifo_inputs_t;
        signal outputs_full_140097944145312: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944145368: core_fifo_inputs_t;
        signal fifo_full_140097944145368: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944145368: core_fifo_inputs_t;
        signal outputs_full_140097944145368: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944145424: core_fifo_inputs_t;
        signal fifo_full_140097944145424: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944145424: core_fifo_inputs_t;
        signal outputs_full_140097944145424: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944145480: core_fifo_inputs_t;
        signal fifo_full_140097944145480: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944145480: core_fifo_inputs_t;
        signal outputs_full_140097944145480: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944145536: core_fifo_inputs_t;
        signal fifo_full_140097944145536: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944145536: core_fifo_inputs_t;
        signal outputs_full_140097944145536: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944145592: core_fifo_inputs_t;
        signal fifo_full_140097944145592: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944145592: core_fifo_inputs_t;
        signal outputs_full_140097944145592: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944145648: core_fifo_inputs_t;
        signal fifo_full_140097944145648: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944145648: core_fifo_inputs_t;
        signal outputs_full_140097944145648: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944145704: core_fifo_inputs_t;
        signal fifo_full_140097944145704: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944145704: core_fifo_inputs_t;
        signal outputs_full_140097944145704: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944145760: core_fifo_inputs_t;
        signal fifo_full_140097944145760: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944145760: core_fifo_inputs_t;
        signal outputs_full_140097944145760: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944145816: core_fifo_inputs_t;
        signal fifo_full_140097944145816: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944145816: core_fifo_inputs_t;
        signal outputs_full_140097944145816: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944145872: core_fifo_inputs_t;
        signal fifo_full_140097944145872: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944145872: core_fifo_inputs_t;
        signal outputs_full_140097944145872: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944154184: core_fifo_inputs_t;
        signal fifo_full_140097944154184: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944154184: core_fifo_inputs_t;
        signal outputs_full_140097944154184: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944154240: core_fifo_inputs_t;
        signal fifo_full_140097944154240: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944154240: core_fifo_inputs_t;
        signal outputs_full_140097944154240: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944154296: core_fifo_inputs_t;
        signal fifo_full_140097944154296: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944154296: core_fifo_inputs_t;
        signal outputs_full_140097944154296: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944154352: core_fifo_inputs_t;
        signal fifo_full_140097944154352: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944154352: core_fifo_inputs_t;
        signal outputs_full_140097944154352: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944154408: core_fifo_inputs_t;
        signal fifo_full_140097944154408: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944154408: core_fifo_inputs_t;
        signal outputs_full_140097944154408: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944154464: core_fifo_inputs_t;
        signal fifo_full_140097944154464: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944154464: core_fifo_inputs_t;
        signal outputs_full_140097944154464: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944154520: core_fifo_inputs_t;
        signal fifo_full_140097944154520: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944154520: core_fifo_inputs_t;
        signal outputs_full_140097944154520: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944154576: core_fifo_inputs_t;
        signal fifo_full_140097944154576: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944154576: core_fifo_inputs_t;
        signal outputs_full_140097944154576: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944154632: core_fifo_inputs_t;
        signal fifo_full_140097944154632: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944154632: core_fifo_inputs_t;
        signal outputs_full_140097944154632: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944154688: core_fifo_inputs_t;
        signal fifo_full_140097944154688: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944154688: core_fifo_inputs_t;
        signal outputs_full_140097944154688: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944154744: core_fifo_inputs_t;
        signal fifo_full_140097944154744: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944154744: core_fifo_inputs_t;
        signal outputs_full_140097944154744: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944154800: core_fifo_inputs_t;
        signal fifo_full_140097944154800: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944154800: core_fifo_inputs_t;
        signal outputs_full_140097944154800: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944154856: core_fifo_inputs_t;
        signal fifo_full_140097944154856: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944154856: core_fifo_inputs_t;
        signal outputs_full_140097944154856: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944154912: core_fifo_inputs_t;
        signal fifo_full_140097944154912: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944154912: core_fifo_inputs_t;
        signal outputs_full_140097944154912: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944154968: core_fifo_inputs_t;
        signal fifo_full_140097944154968: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944154968: core_fifo_inputs_t;
        signal outputs_full_140097944154968: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944155024: core_fifo_inputs_t;
        signal fifo_full_140097944155024: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944155024: core_fifo_inputs_t;
        signal outputs_full_140097944155024: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944155080: core_fifo_inputs_t;
        signal fifo_full_140097944155080: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944155080: core_fifo_inputs_t;
        signal outputs_full_140097944155080: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944155136: core_fifo_inputs_t;
        signal fifo_full_140097944155136: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944155136: core_fifo_inputs_t;
        signal outputs_full_140097944155136: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944155192: core_fifo_inputs_t;
        signal fifo_full_140097944155192: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944155192: core_fifo_inputs_t;
        signal outputs_full_140097944155192: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944155248: core_fifo_inputs_t;
        signal fifo_full_140097944155248: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944155248: core_fifo_inputs_t;
        signal outputs_full_140097944155248: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944155304: core_fifo_inputs_t;
        signal fifo_full_140097944155304: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944155304: core_fifo_inputs_t;
        signal outputs_full_140097944155304: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944155360: core_fifo_inputs_t;
        signal fifo_full_140097944155360: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944155360: core_fifo_inputs_t;
        signal outputs_full_140097944155360: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944155416: core_fifo_inputs_t;
        signal fifo_full_140097944155416: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944155416: core_fifo_inputs_t;
        signal outputs_full_140097944155416: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944155472: core_fifo_inputs_t;
        signal fifo_full_140097944155472: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944155472: core_fifo_inputs_t;
        signal outputs_full_140097944155472: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944155528: core_fifo_inputs_t;
        signal fifo_full_140097944155528: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944155528: core_fifo_inputs_t;
        signal outputs_full_140097944155528: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944155584: core_fifo_inputs_t;
        signal fifo_full_140097944155584: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944155584: core_fifo_inputs_t;
        signal outputs_full_140097944155584: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944155640: core_fifo_inputs_t;
        signal fifo_full_140097944155640: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944155640: core_fifo_inputs_t;
        signal outputs_full_140097944155640: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944155696: core_fifo_inputs_t;
        signal fifo_full_140097944155696: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944155696: core_fifo_inputs_t;
        signal outputs_full_140097944155696: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944155752: core_fifo_inputs_t;
        signal fifo_full_140097944155752: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944155752: core_fifo_inputs_t;
        signal outputs_full_140097944155752: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944155808: core_fifo_inputs_t;
        signal fifo_full_140097944155808: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944155808: core_fifo_inputs_t;
        signal outputs_full_140097944155808: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944155864: core_fifo_inputs_t;
        signal fifo_full_140097944155864: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944155864: core_fifo_inputs_t;
        signal outputs_full_140097944155864: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944155920: core_fifo_inputs_t;
        signal fifo_full_140097944155920: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944155920: core_fifo_inputs_t;
        signal outputs_full_140097944155920: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944155976: core_fifo_inputs_t;
        signal fifo_full_140097944155976: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944155976: core_fifo_inputs_t;
        signal outputs_full_140097944155976: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944156032: core_fifo_inputs_t;
        signal fifo_full_140097944156032: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944156032: core_fifo_inputs_t;
        signal outputs_full_140097944156032: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944156088: core_fifo_inputs_t;
        signal fifo_full_140097944156088: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944156088: core_fifo_inputs_t;
        signal outputs_full_140097944156088: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944156144: core_fifo_inputs_t;
        signal fifo_full_140097944156144: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944156144: core_fifo_inputs_t;
        signal outputs_full_140097944156144: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944156200: core_fifo_inputs_t;
        signal fifo_full_140097944156200: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944156200: core_fifo_inputs_t;
        signal outputs_full_140097944156200: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944156256: core_fifo_inputs_t;
        signal fifo_full_140097944156256: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944156256: core_fifo_inputs_t;
        signal outputs_full_140097944156256: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944156312: core_fifo_inputs_t;
        signal fifo_full_140097944156312: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944156312: core_fifo_inputs_t;
        signal outputs_full_140097944156312: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944156368: core_fifo_inputs_t;
        signal fifo_full_140097944156368: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944156368: core_fifo_inputs_t;
        signal outputs_full_140097944156368: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944156424: core_fifo_inputs_t;
        signal fifo_full_140097944156424: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944156424: core_fifo_inputs_t;
        signal outputs_full_140097944156424: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944156480: core_fifo_inputs_t;
        signal fifo_full_140097944156480: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944156480: core_fifo_inputs_t;
        signal outputs_full_140097944156480: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944156536: core_fifo_inputs_t;
        signal fifo_full_140097944156536: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944156536: core_fifo_inputs_t;
        signal outputs_full_140097944156536: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944156592: core_fifo_inputs_t;
        signal fifo_full_140097944156592: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944156592: core_fifo_inputs_t;
        signal outputs_full_140097944156592: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944156648: core_fifo_inputs_t;
        signal fifo_full_140097944156648: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944156648: core_fifo_inputs_t;
        signal outputs_full_140097944156648: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944156704: core_fifo_inputs_t;
        signal fifo_full_140097944156704: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944156704: core_fifo_inputs_t;
        signal outputs_full_140097944156704: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944156760: core_fifo_inputs_t;
        signal fifo_full_140097944156760: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944156760: core_fifo_inputs_t;
        signal outputs_full_140097944156760: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944156816: core_fifo_inputs_t;
        signal fifo_full_140097944156816: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944156816: core_fifo_inputs_t;
        signal outputs_full_140097944156816: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944156872: core_fifo_inputs_t;
        signal fifo_full_140097944156872: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944156872: core_fifo_inputs_t;
        signal outputs_full_140097944156872: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944156928: core_fifo_inputs_t;
        signal fifo_full_140097944156928: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944156928: core_fifo_inputs_t;
        signal outputs_full_140097944156928: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944156984: core_fifo_inputs_t;
        signal fifo_full_140097944156984: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944156984: core_fifo_inputs_t;
        signal outputs_full_140097944156984: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944157040: core_fifo_inputs_t;
        signal fifo_full_140097944157040: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944157040: core_fifo_inputs_t;
        signal outputs_full_140097944157040: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944157096: core_fifo_inputs_t;
        signal fifo_full_140097944157096: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944157096: core_fifo_inputs_t;
        signal outputs_full_140097944157096: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944157152: core_fifo_inputs_t;
        signal fifo_full_140097944157152: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944157152: core_fifo_inputs_t;
        signal outputs_full_140097944157152: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944157208: core_fifo_inputs_t;
        signal fifo_full_140097944157208: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944157208: core_fifo_inputs_t;
        signal outputs_full_140097944157208: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944157264: core_fifo_inputs_t;
        signal fifo_full_140097944157264: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944157264: core_fifo_inputs_t;
        signal outputs_full_140097944157264: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944157320: core_fifo_inputs_t;
        signal fifo_full_140097944157320: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944157320: core_fifo_inputs_t;
        signal outputs_full_140097944157320: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944157376: core_fifo_inputs_t;
        signal fifo_full_140097944157376: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944157376: core_fifo_inputs_t;
        signal outputs_full_140097944157376: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944157432: core_fifo_inputs_t;
        signal fifo_full_140097944157432: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944157432: core_fifo_inputs_t;
        signal outputs_full_140097944157432: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944157488: core_fifo_inputs_t;
        signal fifo_full_140097944157488: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944157488: core_fifo_inputs_t;
        signal outputs_full_140097944157488: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944157544: core_fifo_inputs_t;
        signal fifo_full_140097944157544: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944157544: core_fifo_inputs_t;
        signal outputs_full_140097944157544: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944157600: core_fifo_inputs_t;
        signal fifo_full_140097944157600: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944157600: core_fifo_inputs_t;
        signal outputs_full_140097944157600: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944157656: core_fifo_inputs_t;
        signal fifo_full_140097944157656: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944157656: core_fifo_inputs_t;
        signal outputs_full_140097944157656: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944157712: core_fifo_inputs_t;
        signal fifo_full_140097944157712: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944157712: core_fifo_inputs_t;
        signal outputs_full_140097944157712: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944157768: core_fifo_inputs_t;
        signal fifo_full_140097944157768: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944157768: core_fifo_inputs_t;
        signal outputs_full_140097944157768: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944157824: core_fifo_inputs_t;
        signal fifo_full_140097944157824: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944157824: core_fifo_inputs_t;
        signal outputs_full_140097944157824: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944157880: core_fifo_inputs_t;
        signal fifo_full_140097944157880: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944157880: core_fifo_inputs_t;
        signal outputs_full_140097944157880: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944157936: core_fifo_inputs_t;
        signal fifo_full_140097944157936: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944157936: core_fifo_inputs_t;
        signal outputs_full_140097944157936: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944157992: core_fifo_inputs_t;
        signal fifo_full_140097944157992: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944157992: core_fifo_inputs_t;
        signal outputs_full_140097944157992: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944158048: core_fifo_inputs_t;
        signal fifo_full_140097944158048: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944158048: core_fifo_inputs_t;
        signal outputs_full_140097944158048: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944158104: core_fifo_inputs_t;
        signal fifo_full_140097944158104: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944158104: core_fifo_inputs_t;
        signal outputs_full_140097944158104: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944158160: core_fifo_inputs_t;
        signal fifo_full_140097944158160: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944158160: core_fifo_inputs_t;
        signal outputs_full_140097944158160: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944166472: core_fifo_inputs_t;
        signal fifo_full_140097944166472: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944166472: core_fifo_inputs_t;
        signal outputs_full_140097944166472: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944166528: core_fifo_inputs_t;
        signal fifo_full_140097944166528: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944166528: core_fifo_inputs_t;
        signal outputs_full_140097944166528: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944166584: core_fifo_inputs_t;
        signal fifo_full_140097944166584: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944166584: core_fifo_inputs_t;
        signal outputs_full_140097944166584: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944166640: core_fifo_inputs_t;
        signal fifo_full_140097944166640: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944166640: core_fifo_inputs_t;
        signal outputs_full_140097944166640: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944166696: core_fifo_inputs_t;
        signal fifo_full_140097944166696: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944166696: core_fifo_inputs_t;
        signal outputs_full_140097944166696: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944166752: core_fifo_inputs_t;
        signal fifo_full_140097944166752: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944166752: core_fifo_inputs_t;
        signal outputs_full_140097944166752: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944166808: core_fifo_inputs_t;
        signal fifo_full_140097944166808: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944166808: core_fifo_inputs_t;
        signal outputs_full_140097944166808: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944166864: core_fifo_inputs_t;
        signal fifo_full_140097944166864: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944166864: core_fifo_inputs_t;
        signal outputs_full_140097944166864: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944166920: core_fifo_inputs_t;
        signal fifo_full_140097944166920: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944166920: core_fifo_inputs_t;
        signal outputs_full_140097944166920: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944166976: core_fifo_inputs_t;
        signal fifo_full_140097944166976: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944166976: core_fifo_inputs_t;
        signal outputs_full_140097944166976: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944167032: core_fifo_inputs_t;
        signal fifo_full_140097944167032: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944167032: core_fifo_inputs_t;
        signal outputs_full_140097944167032: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944167088: core_fifo_inputs_t;
        signal fifo_full_140097944167088: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944167088: core_fifo_inputs_t;
        signal outputs_full_140097944167088: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944167144: core_fifo_inputs_t;
        signal fifo_full_140097944167144: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944167144: core_fifo_inputs_t;
        signal outputs_full_140097944167144: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944167200: core_fifo_inputs_t;
        signal fifo_full_140097944167200: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944167200: core_fifo_inputs_t;
        signal outputs_full_140097944167200: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944167256: core_fifo_inputs_t;
        signal fifo_full_140097944167256: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944167256: core_fifo_inputs_t;
        signal outputs_full_140097944167256: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944167312: core_fifo_inputs_t;
        signal fifo_full_140097944167312: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944167312: core_fifo_inputs_t;
        signal outputs_full_140097944167312: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944167368: core_fifo_inputs_t;
        signal fifo_full_140097944167368: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944167368: core_fifo_inputs_t;
        signal outputs_full_140097944167368: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944167424: core_fifo_inputs_t;
        signal fifo_full_140097944167424: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944167424: core_fifo_inputs_t;
        signal outputs_full_140097944167424: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944167480: core_fifo_inputs_t;
        signal fifo_full_140097944167480: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944167480: core_fifo_inputs_t;
        signal outputs_full_140097944167480: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944167536: core_fifo_inputs_t;
        signal fifo_full_140097944167536: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944167536: core_fifo_inputs_t;
        signal outputs_full_140097944167536: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944167592: core_fifo_inputs_t;
        signal fifo_full_140097944167592: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944167592: core_fifo_inputs_t;
        signal outputs_full_140097944167592: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944167648: core_fifo_inputs_t;
        signal fifo_full_140097944167648: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944167648: core_fifo_inputs_t;
        signal outputs_full_140097944167648: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944167704: core_fifo_inputs_t;
        signal fifo_full_140097944167704: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944167704: core_fifo_inputs_t;
        signal outputs_full_140097944167704: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944167760: core_fifo_inputs_t;
        signal fifo_full_140097944167760: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944167760: core_fifo_inputs_t;
        signal outputs_full_140097944167760: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944167816: core_fifo_inputs_t;
        signal fifo_full_140097944167816: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944167816: core_fifo_inputs_t;
        signal outputs_full_140097944167816: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944167872: core_fifo_inputs_t;
        signal fifo_full_140097944167872: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944167872: core_fifo_inputs_t;
        signal outputs_full_140097944167872: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944167928: core_fifo_inputs_t;
        signal fifo_full_140097944167928: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944167928: core_fifo_inputs_t;
        signal outputs_full_140097944167928: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944167984: core_fifo_inputs_t;
        signal fifo_full_140097944167984: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944167984: core_fifo_inputs_t;
        signal outputs_full_140097944167984: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944168040: core_fifo_inputs_t;
        signal fifo_full_140097944168040: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944168040: core_fifo_inputs_t;
        signal outputs_full_140097944168040: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944168096: core_fifo_inputs_t;
        signal fifo_full_140097944168096: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944168096: core_fifo_inputs_t;
        signal outputs_full_140097944168096: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944168152: core_fifo_inputs_t;
        signal fifo_full_140097944168152: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944168152: core_fifo_inputs_t;
        signal outputs_full_140097944168152: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944168208: core_fifo_inputs_t;
        signal fifo_full_140097944168208: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944168208: core_fifo_inputs_t;
        signal outputs_full_140097944168208: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944168264: core_fifo_inputs_t;
        signal fifo_full_140097944168264: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944168264: core_fifo_inputs_t;
        signal outputs_full_140097944168264: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944168320: core_fifo_inputs_t;
        signal fifo_full_140097944168320: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944168320: core_fifo_inputs_t;
        signal outputs_full_140097944168320: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944168376: core_fifo_inputs_t;
        signal fifo_full_140097944168376: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944168376: core_fifo_inputs_t;
        signal outputs_full_140097944168376: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944168432: core_fifo_inputs_t;
        signal fifo_full_140097944168432: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944168432: core_fifo_inputs_t;
        signal outputs_full_140097944168432: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944168488: core_fifo_inputs_t;
        signal fifo_full_140097944168488: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944168488: core_fifo_inputs_t;
        signal outputs_full_140097944168488: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944168544: core_fifo_inputs_t;
        signal fifo_full_140097944168544: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944168544: core_fifo_inputs_t;
        signal outputs_full_140097944168544: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944168600: core_fifo_inputs_t;
        signal fifo_full_140097944168600: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944168600: core_fifo_inputs_t;
        signal outputs_full_140097944168600: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944168656: core_fifo_inputs_t;
        signal fifo_full_140097944168656: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944168656: core_fifo_inputs_t;
        signal outputs_full_140097944168656: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944168712: core_fifo_inputs_t;
        signal fifo_full_140097944168712: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944168712: core_fifo_inputs_t;
        signal outputs_full_140097944168712: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944168768: core_fifo_inputs_t;
        signal fifo_full_140097944168768: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944168768: core_fifo_inputs_t;
        signal outputs_full_140097944168768: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944168824: core_fifo_inputs_t;
        signal fifo_full_140097944168824: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944168824: core_fifo_inputs_t;
        signal outputs_full_140097944168824: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944168880: core_fifo_inputs_t;
        signal fifo_full_140097944168880: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944168880: core_fifo_inputs_t;
        signal outputs_full_140097944168880: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944168936: core_fifo_inputs_t;
        signal fifo_full_140097944168936: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944168936: core_fifo_inputs_t;
        signal outputs_full_140097944168936: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944168992: core_fifo_inputs_t;
        signal fifo_full_140097944168992: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944168992: core_fifo_inputs_t;
        signal outputs_full_140097944168992: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944169048: core_fifo_inputs_t;
        signal fifo_full_140097944169048: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944169048: core_fifo_inputs_t;
        signal outputs_full_140097944169048: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944169104: core_fifo_inputs_t;
        signal fifo_full_140097944169104: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944169104: core_fifo_inputs_t;
        signal outputs_full_140097944169104: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944169160: core_fifo_inputs_t;
        signal fifo_full_140097944169160: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944169160: core_fifo_inputs_t;
        signal outputs_full_140097944169160: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944169216: core_fifo_inputs_t;
        signal fifo_full_140097944169216: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944169216: core_fifo_inputs_t;
        signal outputs_full_140097944169216: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944169272: core_fifo_inputs_t;
        signal fifo_full_140097944169272: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944169272: core_fifo_inputs_t;
        signal outputs_full_140097944169272: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944169328: core_fifo_inputs_t;
        signal fifo_full_140097944169328: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944169328: core_fifo_inputs_t;
        signal outputs_full_140097944169328: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944169384: core_fifo_inputs_t;
        signal fifo_full_140097944169384: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944169384: core_fifo_inputs_t;
        signal outputs_full_140097944169384: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944169440: core_fifo_inputs_t;
        signal fifo_full_140097944169440: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944169440: core_fifo_inputs_t;
        signal outputs_full_140097944169440: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944169496: core_fifo_inputs_t;
        signal fifo_full_140097944169496: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944169496: core_fifo_inputs_t;
        signal outputs_full_140097944169496: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944169552: core_fifo_inputs_t;
        signal fifo_full_140097944169552: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944169552: core_fifo_inputs_t;
        signal outputs_full_140097944169552: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944169608: core_fifo_inputs_t;
        signal fifo_full_140097944169608: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944169608: core_fifo_inputs_t;
        signal outputs_full_140097944169608: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944169664: core_fifo_inputs_t;
        signal fifo_full_140097944169664: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944169664: core_fifo_inputs_t;
        signal outputs_full_140097944169664: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944169720: core_fifo_inputs_t;
        signal fifo_full_140097944169720: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944169720: core_fifo_inputs_t;
        signal outputs_full_140097944169720: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944169776: core_fifo_inputs_t;
        signal fifo_full_140097944169776: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944169776: core_fifo_inputs_t;
        signal outputs_full_140097944169776: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944169832: core_fifo_inputs_t;
        signal fifo_full_140097944169832: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944169832: core_fifo_inputs_t;
        signal outputs_full_140097944169832: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944169888: core_fifo_inputs_t;
        signal fifo_full_140097944169888: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944169888: core_fifo_inputs_t;
        signal outputs_full_140097944169888: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944169944: core_fifo_inputs_t;
        signal fifo_full_140097944169944: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944169944: core_fifo_inputs_t;
        signal outputs_full_140097944169944: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944170000: core_fifo_inputs_t;
        signal fifo_full_140097944170000: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944170000: core_fifo_inputs_t;
        signal outputs_full_140097944170000: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944170056: core_fifo_inputs_t;
        signal fifo_full_140097944170056: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944170056: core_fifo_inputs_t;
        signal outputs_full_140097944170056: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944170112: core_fifo_inputs_t;
        signal fifo_full_140097944170112: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944170112: core_fifo_inputs_t;
        signal outputs_full_140097944170112: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944170168: core_fifo_inputs_t;
        signal fifo_full_140097944170168: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944170168: core_fifo_inputs_t;
        signal outputs_full_140097944170168: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944170224: core_fifo_inputs_t;
        signal fifo_full_140097944170224: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944170224: core_fifo_inputs_t;
        signal outputs_full_140097944170224: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944170280: core_fifo_inputs_t;
        signal fifo_full_140097944170280: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944170280: core_fifo_inputs_t;
        signal outputs_full_140097944170280: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944170336: core_fifo_inputs_t;
        signal fifo_full_140097944170336: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944170336: core_fifo_inputs_t;
        signal outputs_full_140097944170336: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944170392: core_fifo_inputs_t;
        signal fifo_full_140097944170392: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944170392: core_fifo_inputs_t;
        signal outputs_full_140097944170392: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097944170448: core_fifo_inputs_t;
        signal fifo_full_140097944170448: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097944170448: core_fifo_inputs_t;
        signal outputs_full_140097944170448: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941516360: core_fifo_inputs_t;
        signal fifo_full_140097941516360: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941516360: core_fifo_inputs_t;
        signal outputs_full_140097941516360: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941516416: core_fifo_inputs_t;
        signal fifo_full_140097941516416: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941516416: core_fifo_inputs_t;
        signal outputs_full_140097941516416: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941516472: core_fifo_inputs_t;
        signal fifo_full_140097941516472: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941516472: core_fifo_inputs_t;
        signal outputs_full_140097941516472: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941516528: core_fifo_inputs_t;
        signal fifo_full_140097941516528: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941516528: core_fifo_inputs_t;
        signal outputs_full_140097941516528: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941516584: core_fifo_inputs_t;
        signal fifo_full_140097941516584: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941516584: core_fifo_inputs_t;
        signal outputs_full_140097941516584: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941516640: core_fifo_inputs_t;
        signal fifo_full_140097941516640: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941516640: core_fifo_inputs_t;
        signal outputs_full_140097941516640: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941516696: core_fifo_inputs_t;
        signal fifo_full_140097941516696: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941516696: core_fifo_inputs_t;
        signal outputs_full_140097941516696: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941516752: core_fifo_inputs_t;
        signal fifo_full_140097941516752: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941516752: core_fifo_inputs_t;
        signal outputs_full_140097941516752: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941516808: core_fifo_inputs_t;
        signal fifo_full_140097941516808: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941516808: core_fifo_inputs_t;
        signal outputs_full_140097941516808: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941516864: core_fifo_inputs_t;
        signal fifo_full_140097941516864: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941516864: core_fifo_inputs_t;
        signal outputs_full_140097941516864: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941516920: core_fifo_inputs_t;
        signal fifo_full_140097941516920: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941516920: core_fifo_inputs_t;
        signal outputs_full_140097941516920: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941516976: core_fifo_inputs_t;
        signal fifo_full_140097941516976: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941516976: core_fifo_inputs_t;
        signal outputs_full_140097941516976: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941517032: core_fifo_inputs_t;
        signal fifo_full_140097941517032: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941517032: core_fifo_inputs_t;
        signal outputs_full_140097941517032: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941517088: core_fifo_inputs_t;
        signal fifo_full_140097941517088: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941517088: core_fifo_inputs_t;
        signal outputs_full_140097941517088: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941517144: core_fifo_inputs_t;
        signal fifo_full_140097941517144: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941517144: core_fifo_inputs_t;
        signal outputs_full_140097941517144: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941517200: core_fifo_inputs_t;
        signal fifo_full_140097941517200: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941517200: core_fifo_inputs_t;
        signal outputs_full_140097941517200: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941517256: core_fifo_inputs_t;
        signal fifo_full_140097941517256: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941517256: core_fifo_inputs_t;
        signal outputs_full_140097941517256: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941517312: core_fifo_inputs_t;
        signal fifo_full_140097941517312: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941517312: core_fifo_inputs_t;
        signal outputs_full_140097941517312: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941517368: core_fifo_inputs_t;
        signal fifo_full_140097941517368: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941517368: core_fifo_inputs_t;
        signal outputs_full_140097941517368: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941517424: core_fifo_inputs_t;
        signal fifo_full_140097941517424: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941517424: core_fifo_inputs_t;
        signal outputs_full_140097941517424: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941517480: core_fifo_inputs_t;
        signal fifo_full_140097941517480: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941517480: core_fifo_inputs_t;
        signal outputs_full_140097941517480: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941517536: core_fifo_inputs_t;
        signal fifo_full_140097941517536: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941517536: core_fifo_inputs_t;
        signal outputs_full_140097941517536: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941517592: core_fifo_inputs_t;
        signal fifo_full_140097941517592: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941517592: core_fifo_inputs_t;
        signal outputs_full_140097941517592: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941517648: core_fifo_inputs_t;
        signal fifo_full_140097941517648: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941517648: core_fifo_inputs_t;
        signal outputs_full_140097941517648: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941517704: core_fifo_inputs_t;
        signal fifo_full_140097941517704: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941517704: core_fifo_inputs_t;
        signal outputs_full_140097941517704: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941517760: core_fifo_inputs_t;
        signal fifo_full_140097941517760: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941517760: core_fifo_inputs_t;
        signal outputs_full_140097941517760: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941517816: core_fifo_inputs_t;
        signal fifo_full_140097941517816: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941517816: core_fifo_inputs_t;
        signal outputs_full_140097941517816: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941517872: core_fifo_inputs_t;
        signal fifo_full_140097941517872: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941517872: core_fifo_inputs_t;
        signal outputs_full_140097941517872: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941517928: core_fifo_inputs_t;
        signal fifo_full_140097941517928: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941517928: core_fifo_inputs_t;
        signal outputs_full_140097941517928: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941517984: core_fifo_inputs_t;
        signal fifo_full_140097941517984: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941517984: core_fifo_inputs_t;
        signal outputs_full_140097941517984: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941518040: core_fifo_inputs_t;
        signal fifo_full_140097941518040: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941518040: core_fifo_inputs_t;
        signal outputs_full_140097941518040: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941518096: core_fifo_inputs_t;
        signal fifo_full_140097941518096: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941518096: core_fifo_inputs_t;
        signal outputs_full_140097941518096: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941518152: core_fifo_inputs_t;
        signal fifo_full_140097941518152: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941518152: core_fifo_inputs_t;
        signal outputs_full_140097941518152: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941518208: core_fifo_inputs_t;
        signal fifo_full_140097941518208: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941518208: core_fifo_inputs_t;
        signal outputs_full_140097941518208: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941518264: core_fifo_inputs_t;
        signal fifo_full_140097941518264: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941518264: core_fifo_inputs_t;
        signal outputs_full_140097941518264: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941518320: core_fifo_inputs_t;
        signal fifo_full_140097941518320: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941518320: core_fifo_inputs_t;
        signal outputs_full_140097941518320: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941518376: core_fifo_inputs_t;
        signal fifo_full_140097941518376: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941518376: core_fifo_inputs_t;
        signal outputs_full_140097941518376: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941518432: core_fifo_inputs_t;
        signal fifo_full_140097941518432: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941518432: core_fifo_inputs_t;
        signal outputs_full_140097941518432: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941518488: core_fifo_inputs_t;
        signal fifo_full_140097941518488: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941518488: core_fifo_inputs_t;
        signal outputs_full_140097941518488: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941518544: core_fifo_inputs_t;
        signal fifo_full_140097941518544: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941518544: core_fifo_inputs_t;
        signal outputs_full_140097941518544: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941518600: core_fifo_inputs_t;
        signal fifo_full_140097941518600: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941518600: core_fifo_inputs_t;
        signal outputs_full_140097941518600: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941518656: core_fifo_inputs_t;
        signal fifo_full_140097941518656: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941518656: core_fifo_inputs_t;
        signal outputs_full_140097941518656: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941518712: core_fifo_inputs_t;
        signal fifo_full_140097941518712: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941518712: core_fifo_inputs_t;
        signal outputs_full_140097941518712: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941518768: core_fifo_inputs_t;
        signal fifo_full_140097941518768: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941518768: core_fifo_inputs_t;
        signal outputs_full_140097941518768: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941518824: core_fifo_inputs_t;
        signal fifo_full_140097941518824: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941518824: core_fifo_inputs_t;
        signal outputs_full_140097941518824: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941518880: core_fifo_inputs_t;
        signal fifo_full_140097941518880: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941518880: core_fifo_inputs_t;
        signal outputs_full_140097941518880: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941518936: core_fifo_inputs_t;
        signal fifo_full_140097941518936: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941518936: core_fifo_inputs_t;
        signal outputs_full_140097941518936: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941518992: core_fifo_inputs_t;
        signal fifo_full_140097941518992: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941518992: core_fifo_inputs_t;
        signal outputs_full_140097941518992: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941519048: core_fifo_inputs_t;
        signal fifo_full_140097941519048: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941519048: core_fifo_inputs_t;
        signal outputs_full_140097941519048: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941519104: core_fifo_inputs_t;
        signal fifo_full_140097941519104: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941519104: core_fifo_inputs_t;
        signal outputs_full_140097941519104: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941519160: core_fifo_inputs_t;
        signal fifo_full_140097941519160: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941519160: core_fifo_inputs_t;
        signal outputs_full_140097941519160: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941519216: core_fifo_inputs_t;
        signal fifo_full_140097941519216: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941519216: core_fifo_inputs_t;
        signal outputs_full_140097941519216: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941519272: core_fifo_inputs_t;
        signal fifo_full_140097941519272: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941519272: core_fifo_inputs_t;
        signal outputs_full_140097941519272: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941519328: core_fifo_inputs_t;
        signal fifo_full_140097941519328: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941519328: core_fifo_inputs_t;
        signal outputs_full_140097941519328: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941519384: core_fifo_inputs_t;
        signal fifo_full_140097941519384: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941519384: core_fifo_inputs_t;
        signal outputs_full_140097941519384: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941519440: core_fifo_inputs_t;
        signal fifo_full_140097941519440: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941519440: core_fifo_inputs_t;
        signal outputs_full_140097941519440: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941519496: core_fifo_inputs_t;
        signal fifo_full_140097941519496: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941519496: core_fifo_inputs_t;
        signal outputs_full_140097941519496: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941519552: core_fifo_inputs_t;
        signal fifo_full_140097941519552: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941519552: core_fifo_inputs_t;
        signal outputs_full_140097941519552: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941519608: core_fifo_inputs_t;
        signal fifo_full_140097941519608: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941519608: core_fifo_inputs_t;
        signal outputs_full_140097941519608: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941519664: core_fifo_inputs_t;
        signal fifo_full_140097941519664: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941519664: core_fifo_inputs_t;
        signal outputs_full_140097941519664: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941519720: core_fifo_inputs_t;
        signal fifo_full_140097941519720: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941519720: core_fifo_inputs_t;
        signal outputs_full_140097941519720: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941519776: core_fifo_inputs_t;
        signal fifo_full_140097941519776: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941519776: core_fifo_inputs_t;
        signal outputs_full_140097941519776: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941519832: core_fifo_inputs_t;
        signal fifo_full_140097941519832: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941519832: core_fifo_inputs_t;
        signal outputs_full_140097941519832: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941519888: core_fifo_inputs_t;
        signal fifo_full_140097941519888: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941519888: core_fifo_inputs_t;
        signal outputs_full_140097941519888: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941519944: core_fifo_inputs_t;
        signal fifo_full_140097941519944: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941519944: core_fifo_inputs_t;
        signal outputs_full_140097941519944: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941520000: core_fifo_inputs_t;
        signal fifo_full_140097941520000: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941520000: core_fifo_inputs_t;
        signal outputs_full_140097941520000: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941520056: core_fifo_inputs_t;
        signal fifo_full_140097941520056: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941520056: core_fifo_inputs_t;
        signal outputs_full_140097941520056: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941520112: core_fifo_inputs_t;
        signal fifo_full_140097941520112: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941520112: core_fifo_inputs_t;
        signal outputs_full_140097941520112: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941520168: core_fifo_inputs_t;
        signal fifo_full_140097941520168: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941520168: core_fifo_inputs_t;
        signal outputs_full_140097941520168: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941520224: core_fifo_inputs_t;
        signal fifo_full_140097941520224: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941520224: core_fifo_inputs_t;
        signal outputs_full_140097941520224: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941520280: core_fifo_inputs_t;
        signal fifo_full_140097941520280: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941520280: core_fifo_inputs_t;
        signal outputs_full_140097941520280: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941520336: core_fifo_inputs_t;
        signal fifo_full_140097941520336: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941520336: core_fifo_inputs_t;
        signal outputs_full_140097941520336: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941528648: core_fifo_inputs_t;
        signal fifo_full_140097941528648: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941528648: core_fifo_inputs_t;
        signal outputs_full_140097941528648: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941528704: core_fifo_inputs_t;
        signal fifo_full_140097941528704: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941528704: core_fifo_inputs_t;
        signal outputs_full_140097941528704: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941528760: core_fifo_inputs_t;
        signal fifo_full_140097941528760: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941528760: core_fifo_inputs_t;
        signal outputs_full_140097941528760: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941528816: core_fifo_inputs_t;
        signal fifo_full_140097941528816: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941528816: core_fifo_inputs_t;
        signal outputs_full_140097941528816: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941528872: core_fifo_inputs_t;
        signal fifo_full_140097941528872: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941528872: core_fifo_inputs_t;
        signal outputs_full_140097941528872: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941528928: core_fifo_inputs_t;
        signal fifo_full_140097941528928: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941528928: core_fifo_inputs_t;
        signal outputs_full_140097941528928: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941528984: core_fifo_inputs_t;
        signal fifo_full_140097941528984: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941528984: core_fifo_inputs_t;
        signal outputs_full_140097941528984: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941529040: core_fifo_inputs_t;
        signal fifo_full_140097941529040: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941529040: core_fifo_inputs_t;
        signal outputs_full_140097941529040: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941529096: core_fifo_inputs_t;
        signal fifo_full_140097941529096: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941529096: core_fifo_inputs_t;
        signal outputs_full_140097941529096: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941529152: core_fifo_inputs_t;
        signal fifo_full_140097941529152: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941529152: core_fifo_inputs_t;
        signal outputs_full_140097941529152: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941529208: core_fifo_inputs_t;
        signal fifo_full_140097941529208: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941529208: core_fifo_inputs_t;
        signal outputs_full_140097941529208: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941529264: core_fifo_inputs_t;
        signal fifo_full_140097941529264: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941529264: core_fifo_inputs_t;
        signal outputs_full_140097941529264: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941529320: core_fifo_inputs_t;
        signal fifo_full_140097941529320: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941529320: core_fifo_inputs_t;
        signal outputs_full_140097941529320: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941529376: core_fifo_inputs_t;
        signal fifo_full_140097941529376: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941529376: core_fifo_inputs_t;
        signal outputs_full_140097941529376: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941529432: core_fifo_inputs_t;
        signal fifo_full_140097941529432: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941529432: core_fifo_inputs_t;
        signal outputs_full_140097941529432: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941529488: core_fifo_inputs_t;
        signal fifo_full_140097941529488: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941529488: core_fifo_inputs_t;
        signal outputs_full_140097941529488: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941529544: core_fifo_inputs_t;
        signal fifo_full_140097941529544: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941529544: core_fifo_inputs_t;
        signal outputs_full_140097941529544: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941529600: core_fifo_inputs_t;
        signal fifo_full_140097941529600: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941529600: core_fifo_inputs_t;
        signal outputs_full_140097941529600: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941529656: core_fifo_inputs_t;
        signal fifo_full_140097941529656: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941529656: core_fifo_inputs_t;
        signal outputs_full_140097941529656: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941529712: core_fifo_inputs_t;
        signal fifo_full_140097941529712: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941529712: core_fifo_inputs_t;
        signal outputs_full_140097941529712: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941529768: core_fifo_inputs_t;
        signal fifo_full_140097941529768: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941529768: core_fifo_inputs_t;
        signal outputs_full_140097941529768: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941529824: core_fifo_inputs_t;
        signal fifo_full_140097941529824: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941529824: core_fifo_inputs_t;
        signal outputs_full_140097941529824: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941529880: core_fifo_inputs_t;
        signal fifo_full_140097941529880: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941529880: core_fifo_inputs_t;
        signal outputs_full_140097941529880: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941529936: core_fifo_inputs_t;
        signal fifo_full_140097941529936: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941529936: core_fifo_inputs_t;
        signal outputs_full_140097941529936: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941529992: core_fifo_inputs_t;
        signal fifo_full_140097941529992: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941529992: core_fifo_inputs_t;
        signal outputs_full_140097941529992: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941530048: core_fifo_inputs_t;
        signal fifo_full_140097941530048: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941530048: core_fifo_inputs_t;
        signal outputs_full_140097941530048: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941530104: core_fifo_inputs_t;
        signal fifo_full_140097941530104: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941530104: core_fifo_inputs_t;
        signal outputs_full_140097941530104: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941530160: core_fifo_inputs_t;
        signal fifo_full_140097941530160: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941530160: core_fifo_inputs_t;
        signal outputs_full_140097941530160: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941530216: core_fifo_inputs_t;
        signal fifo_full_140097941530216: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941530216: core_fifo_inputs_t;
        signal outputs_full_140097941530216: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941530272: core_fifo_inputs_t;
        signal fifo_full_140097941530272: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941530272: core_fifo_inputs_t;
        signal outputs_full_140097941530272: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941530328: core_fifo_inputs_t;
        signal fifo_full_140097941530328: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941530328: core_fifo_inputs_t;
        signal outputs_full_140097941530328: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941530384: core_fifo_inputs_t;
        signal fifo_full_140097941530384: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941530384: core_fifo_inputs_t;
        signal outputs_full_140097941530384: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941530440: core_fifo_inputs_t;
        signal fifo_full_140097941530440: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941530440: core_fifo_inputs_t;
        signal outputs_full_140097941530440: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941530496: core_fifo_inputs_t;
        signal fifo_full_140097941530496: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941530496: core_fifo_inputs_t;
        signal outputs_full_140097941530496: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941530552: core_fifo_inputs_t;
        signal fifo_full_140097941530552: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941530552: core_fifo_inputs_t;
        signal outputs_full_140097941530552: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941530608: core_fifo_inputs_t;
        signal fifo_full_140097941530608: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941530608: core_fifo_inputs_t;
        signal outputs_full_140097941530608: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941530664: core_fifo_inputs_t;
        signal fifo_full_140097941530664: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941530664: core_fifo_inputs_t;
        signal outputs_full_140097941530664: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941530720: core_fifo_inputs_t;
        signal fifo_full_140097941530720: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941530720: core_fifo_inputs_t;
        signal outputs_full_140097941530720: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941530776: core_fifo_inputs_t;
        signal fifo_full_140097941530776: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941530776: core_fifo_inputs_t;
        signal outputs_full_140097941530776: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941530832: core_fifo_inputs_t;
        signal fifo_full_140097941530832: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941530832: core_fifo_inputs_t;
        signal outputs_full_140097941530832: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941530888: core_fifo_inputs_t;
        signal fifo_full_140097941530888: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941530888: core_fifo_inputs_t;
        signal outputs_full_140097941530888: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941530944: core_fifo_inputs_t;
        signal fifo_full_140097941530944: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941530944: core_fifo_inputs_t;
        signal outputs_full_140097941530944: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941531000: core_fifo_inputs_t;
        signal fifo_full_140097941531000: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941531000: core_fifo_inputs_t;
        signal outputs_full_140097941531000: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941531056: core_fifo_inputs_t;
        signal fifo_full_140097941531056: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941531056: core_fifo_inputs_t;
        signal outputs_full_140097941531056: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941531112: core_fifo_inputs_t;
        signal fifo_full_140097941531112: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941531112: core_fifo_inputs_t;
        signal outputs_full_140097941531112: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941531168: core_fifo_inputs_t;
        signal fifo_full_140097941531168: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941531168: core_fifo_inputs_t;
        signal outputs_full_140097941531168: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941531224: core_fifo_inputs_t;
        signal fifo_full_140097941531224: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941531224: core_fifo_inputs_t;
        signal outputs_full_140097941531224: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941531280: core_fifo_inputs_t;
        signal fifo_full_140097941531280: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941531280: core_fifo_inputs_t;
        signal outputs_full_140097941531280: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941531336: core_fifo_inputs_t;
        signal fifo_full_140097941531336: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941531336: core_fifo_inputs_t;
        signal outputs_full_140097941531336: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941531392: core_fifo_inputs_t;
        signal fifo_full_140097941531392: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941531392: core_fifo_inputs_t;
        signal outputs_full_140097941531392: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941531448: core_fifo_inputs_t;
        signal fifo_full_140097941531448: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941531448: core_fifo_inputs_t;
        signal outputs_full_140097941531448: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941531504: core_fifo_inputs_t;
        signal fifo_full_140097941531504: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941531504: core_fifo_inputs_t;
        signal outputs_full_140097941531504: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941531560: core_fifo_inputs_t;
        signal fifo_full_140097941531560: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941531560: core_fifo_inputs_t;
        signal outputs_full_140097941531560: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941531616: core_fifo_inputs_t;
        signal fifo_full_140097941531616: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941531616: core_fifo_inputs_t;
        signal outputs_full_140097941531616: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941531672: core_fifo_inputs_t;
        signal fifo_full_140097941531672: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941531672: core_fifo_inputs_t;
        signal outputs_full_140097941531672: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941531728: core_fifo_inputs_t;
        signal fifo_full_140097941531728: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941531728: core_fifo_inputs_t;
        signal outputs_full_140097941531728: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941531784: core_fifo_inputs_t;
        signal fifo_full_140097941531784: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941531784: core_fifo_inputs_t;
        signal outputs_full_140097941531784: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941531840: core_fifo_inputs_t;
        signal fifo_full_140097941531840: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941531840: core_fifo_inputs_t;
        signal outputs_full_140097941531840: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941531896: core_fifo_inputs_t;
        signal fifo_full_140097941531896: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941531896: core_fifo_inputs_t;
        signal outputs_full_140097941531896: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941531952: core_fifo_inputs_t;
        signal fifo_full_140097941531952: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941531952: core_fifo_inputs_t;
        signal outputs_full_140097941531952: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941532008: core_fifo_inputs_t;
        signal fifo_full_140097941532008: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941532008: core_fifo_inputs_t;
        signal outputs_full_140097941532008: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941532064: core_fifo_inputs_t;
        signal fifo_full_140097941532064: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941532064: core_fifo_inputs_t;
        signal outputs_full_140097941532064: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941532120: core_fifo_inputs_t;
        signal fifo_full_140097941532120: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941532120: core_fifo_inputs_t;
        signal outputs_full_140097941532120: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941532176: core_fifo_inputs_t;
        signal fifo_full_140097941532176: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941532176: core_fifo_inputs_t;
        signal outputs_full_140097941532176: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941532232: core_fifo_inputs_t;
        signal fifo_full_140097941532232: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941532232: core_fifo_inputs_t;
        signal outputs_full_140097941532232: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941532288: core_fifo_inputs_t;
        signal fifo_full_140097941532288: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941532288: core_fifo_inputs_t;
        signal outputs_full_140097941532288: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941532344: core_fifo_inputs_t;
        signal fifo_full_140097941532344: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941532344: core_fifo_inputs_t;
        signal outputs_full_140097941532344: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941532400: core_fifo_inputs_t;
        signal fifo_full_140097941532400: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941532400: core_fifo_inputs_t;
        signal outputs_full_140097941532400: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941532456: core_fifo_inputs_t;
        signal fifo_full_140097941532456: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941532456: core_fifo_inputs_t;
        signal outputs_full_140097941532456: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941532512: core_fifo_inputs_t;
        signal fifo_full_140097941532512: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941532512: core_fifo_inputs_t;
        signal outputs_full_140097941532512: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941532568: core_fifo_inputs_t;
        signal fifo_full_140097941532568: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941532568: core_fifo_inputs_t;
        signal outputs_full_140097941532568: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941532624: core_fifo_inputs_t;
        signal fifo_full_140097941532624: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941532624: core_fifo_inputs_t;
        signal outputs_full_140097941532624: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941540936: core_fifo_inputs_t;
        signal fifo_full_140097941540936: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941540936: core_fifo_inputs_t;
        signal outputs_full_140097941540936: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941540992: core_fifo_inputs_t;
        signal fifo_full_140097941540992: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941540992: core_fifo_inputs_t;
        signal outputs_full_140097941540992: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941541048: core_fifo_inputs_t;
        signal fifo_full_140097941541048: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941541048: core_fifo_inputs_t;
        signal outputs_full_140097941541048: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941541104: core_fifo_inputs_t;
        signal fifo_full_140097941541104: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941541104: core_fifo_inputs_t;
        signal outputs_full_140097941541104: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941541160: core_fifo_inputs_t;
        signal fifo_full_140097941541160: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941541160: core_fifo_inputs_t;
        signal outputs_full_140097941541160: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941541216: core_fifo_inputs_t;
        signal fifo_full_140097941541216: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941541216: core_fifo_inputs_t;
        signal outputs_full_140097941541216: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941541272: core_fifo_inputs_t;
        signal fifo_full_140097941541272: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941541272: core_fifo_inputs_t;
        signal outputs_full_140097941541272: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941541328: core_fifo_inputs_t;
        signal fifo_full_140097941541328: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941541328: core_fifo_inputs_t;
        signal outputs_full_140097941541328: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941541384: core_fifo_inputs_t;
        signal fifo_full_140097941541384: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941541384: core_fifo_inputs_t;
        signal outputs_full_140097941541384: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941541440: core_fifo_inputs_t;
        signal fifo_full_140097941541440: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941541440: core_fifo_inputs_t;
        signal outputs_full_140097941541440: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941541496: core_fifo_inputs_t;
        signal fifo_full_140097941541496: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941541496: core_fifo_inputs_t;
        signal outputs_full_140097941541496: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941541552: core_fifo_inputs_t;
        signal fifo_full_140097941541552: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941541552: core_fifo_inputs_t;
        signal outputs_full_140097941541552: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941541608: core_fifo_inputs_t;
        signal fifo_full_140097941541608: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941541608: core_fifo_inputs_t;
        signal outputs_full_140097941541608: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941541664: core_fifo_inputs_t;
        signal fifo_full_140097941541664: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941541664: core_fifo_inputs_t;
        signal outputs_full_140097941541664: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941541720: core_fifo_inputs_t;
        signal fifo_full_140097941541720: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941541720: core_fifo_inputs_t;
        signal outputs_full_140097941541720: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941541776: core_fifo_inputs_t;
        signal fifo_full_140097941541776: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941541776: core_fifo_inputs_t;
        signal outputs_full_140097941541776: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941541832: core_fifo_inputs_t;
        signal fifo_full_140097941541832: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941541832: core_fifo_inputs_t;
        signal outputs_full_140097941541832: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941541888: core_fifo_inputs_t;
        signal fifo_full_140097941541888: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941541888: core_fifo_inputs_t;
        signal outputs_full_140097941541888: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941541944: core_fifo_inputs_t;
        signal fifo_full_140097941541944: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941541944: core_fifo_inputs_t;
        signal outputs_full_140097941541944: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941542000: core_fifo_inputs_t;
        signal fifo_full_140097941542000: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941542000: core_fifo_inputs_t;
        signal outputs_full_140097941542000: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941542056: core_fifo_inputs_t;
        signal fifo_full_140097941542056: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941542056: core_fifo_inputs_t;
        signal outputs_full_140097941542056: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941542112: core_fifo_inputs_t;
        signal fifo_full_140097941542112: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941542112: core_fifo_inputs_t;
        signal outputs_full_140097941542112: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941542168: core_fifo_inputs_t;
        signal fifo_full_140097941542168: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941542168: core_fifo_inputs_t;
        signal outputs_full_140097941542168: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941542224: core_fifo_inputs_t;
        signal fifo_full_140097941542224: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941542224: core_fifo_inputs_t;
        signal outputs_full_140097941542224: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941542280: core_fifo_inputs_t;
        signal fifo_full_140097941542280: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941542280: core_fifo_inputs_t;
        signal outputs_full_140097941542280: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941542336: core_fifo_inputs_t;
        signal fifo_full_140097941542336: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941542336: core_fifo_inputs_t;
        signal outputs_full_140097941542336: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941542392: core_fifo_inputs_t;
        signal fifo_full_140097941542392: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941542392: core_fifo_inputs_t;
        signal outputs_full_140097941542392: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941542448: core_fifo_inputs_t;
        signal fifo_full_140097941542448: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941542448: core_fifo_inputs_t;
        signal outputs_full_140097941542448: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941542504: core_fifo_inputs_t;
        signal fifo_full_140097941542504: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941542504: core_fifo_inputs_t;
        signal outputs_full_140097941542504: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941542560: core_fifo_inputs_t;
        signal fifo_full_140097941542560: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941542560: core_fifo_inputs_t;
        signal outputs_full_140097941542560: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941542616: core_fifo_inputs_t;
        signal fifo_full_140097941542616: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941542616: core_fifo_inputs_t;
        signal outputs_full_140097941542616: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941542672: core_fifo_inputs_t;
        signal fifo_full_140097941542672: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941542672: core_fifo_inputs_t;
        signal outputs_full_140097941542672: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941542728: core_fifo_inputs_t;
        signal fifo_full_140097941542728: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941542728: core_fifo_inputs_t;
        signal outputs_full_140097941542728: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941542784: core_fifo_inputs_t;
        signal fifo_full_140097941542784: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941542784: core_fifo_inputs_t;
        signal outputs_full_140097941542784: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941542840: core_fifo_inputs_t;
        signal fifo_full_140097941542840: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941542840: core_fifo_inputs_t;
        signal outputs_full_140097941542840: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941542896: core_fifo_inputs_t;
        signal fifo_full_140097941542896: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941542896: core_fifo_inputs_t;
        signal outputs_full_140097941542896: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941542952: core_fifo_inputs_t;
        signal fifo_full_140097941542952: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941542952: core_fifo_inputs_t;
        signal outputs_full_140097941542952: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941543008: core_fifo_inputs_t;
        signal fifo_full_140097941543008: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941543008: core_fifo_inputs_t;
        signal outputs_full_140097941543008: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941543064: core_fifo_inputs_t;
        signal fifo_full_140097941543064: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941543064: core_fifo_inputs_t;
        signal outputs_full_140097941543064: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941543120: core_fifo_inputs_t;
        signal fifo_full_140097941543120: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941543120: core_fifo_inputs_t;
        signal outputs_full_140097941543120: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941543176: core_fifo_inputs_t;
        signal fifo_full_140097941543176: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941543176: core_fifo_inputs_t;
        signal outputs_full_140097941543176: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941543232: core_fifo_inputs_t;
        signal fifo_full_140097941543232: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941543232: core_fifo_inputs_t;
        signal outputs_full_140097941543232: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941543288: core_fifo_inputs_t;
        signal fifo_full_140097941543288: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941543288: core_fifo_inputs_t;
        signal outputs_full_140097941543288: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941543344: core_fifo_inputs_t;
        signal fifo_full_140097941543344: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941543344: core_fifo_inputs_t;
        signal outputs_full_140097941543344: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941543400: core_fifo_inputs_t;
        signal fifo_full_140097941543400: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941543400: core_fifo_inputs_t;
        signal outputs_full_140097941543400: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941543456: core_fifo_inputs_t;
        signal fifo_full_140097941543456: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941543456: core_fifo_inputs_t;
        signal outputs_full_140097941543456: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941543512: core_fifo_inputs_t;
        signal fifo_full_140097941543512: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941543512: core_fifo_inputs_t;
        signal outputs_full_140097941543512: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941543568: core_fifo_inputs_t;
        signal fifo_full_140097941543568: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941543568: core_fifo_inputs_t;
        signal outputs_full_140097941543568: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941543624: core_fifo_inputs_t;
        signal fifo_full_140097941543624: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941543624: core_fifo_inputs_t;
        signal outputs_full_140097941543624: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941543680: core_fifo_inputs_t;
        signal fifo_full_140097941543680: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941543680: core_fifo_inputs_t;
        signal outputs_full_140097941543680: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941543736: core_fifo_inputs_t;
        signal fifo_full_140097941543736: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941543736: core_fifo_inputs_t;
        signal outputs_full_140097941543736: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941543792: core_fifo_inputs_t;
        signal fifo_full_140097941543792: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941543792: core_fifo_inputs_t;
        signal outputs_full_140097941543792: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941543848: core_fifo_inputs_t;
        signal fifo_full_140097941543848: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941543848: core_fifo_inputs_t;
        signal outputs_full_140097941543848: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941543904: core_fifo_inputs_t;
        signal fifo_full_140097941543904: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941543904: core_fifo_inputs_t;
        signal outputs_full_140097941543904: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941543960: core_fifo_inputs_t;
        signal fifo_full_140097941543960: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941543960: core_fifo_inputs_t;
        signal outputs_full_140097941543960: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941544016: core_fifo_inputs_t;
        signal fifo_full_140097941544016: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941544016: core_fifo_inputs_t;
        signal outputs_full_140097941544016: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941544072: core_fifo_inputs_t;
        signal fifo_full_140097941544072: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941544072: core_fifo_inputs_t;
        signal outputs_full_140097941544072: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941544128: core_fifo_inputs_t;
        signal fifo_full_140097941544128: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941544128: core_fifo_inputs_t;
        signal outputs_full_140097941544128: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941544184: core_fifo_inputs_t;
        signal fifo_full_140097941544184: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941544184: core_fifo_inputs_t;
        signal outputs_full_140097941544184: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941544240: core_fifo_inputs_t;
        signal fifo_full_140097941544240: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941544240: core_fifo_inputs_t;
        signal outputs_full_140097941544240: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941544296: core_fifo_inputs_t;
        signal fifo_full_140097941544296: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941544296: core_fifo_inputs_t;
        signal outputs_full_140097941544296: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941544352: core_fifo_inputs_t;
        signal fifo_full_140097941544352: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941544352: core_fifo_inputs_t;
        signal outputs_full_140097941544352: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941544408: core_fifo_inputs_t;
        signal fifo_full_140097941544408: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941544408: core_fifo_inputs_t;
        signal outputs_full_140097941544408: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941544464: core_fifo_inputs_t;
        signal fifo_full_140097941544464: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941544464: core_fifo_inputs_t;
        signal outputs_full_140097941544464: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941544520: core_fifo_inputs_t;
        signal fifo_full_140097941544520: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941544520: core_fifo_inputs_t;
        signal outputs_full_140097941544520: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941544576: core_fifo_inputs_t;
        signal fifo_full_140097941544576: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941544576: core_fifo_inputs_t;
        signal outputs_full_140097941544576: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941544632: core_fifo_inputs_t;
        signal fifo_full_140097941544632: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941544632: core_fifo_inputs_t;
        signal outputs_full_140097941544632: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941544688: core_fifo_inputs_t;
        signal fifo_full_140097941544688: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941544688: core_fifo_inputs_t;
        signal outputs_full_140097941544688: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941544744: core_fifo_inputs_t;
        signal fifo_full_140097941544744: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941544744: core_fifo_inputs_t;
        signal outputs_full_140097941544744: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941544800: core_fifo_inputs_t;
        signal fifo_full_140097941544800: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941544800: core_fifo_inputs_t;
        signal outputs_full_140097941544800: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941544856: core_fifo_inputs_t;
        signal fifo_full_140097941544856: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941544856: core_fifo_inputs_t;
        signal outputs_full_140097941544856: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941544912: core_fifo_inputs_t;
        signal fifo_full_140097941544912: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941544912: core_fifo_inputs_t;
        signal outputs_full_140097941544912: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941553224: core_fifo_inputs_t;
        signal fifo_full_140097941553224: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941553224: core_fifo_inputs_t;
        signal outputs_full_140097941553224: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941553280: core_fifo_inputs_t;
        signal fifo_full_140097941553280: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941553280: core_fifo_inputs_t;
        signal outputs_full_140097941553280: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941553336: core_fifo_inputs_t;
        signal fifo_full_140097941553336: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941553336: core_fifo_inputs_t;
        signal outputs_full_140097941553336: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941553392: core_fifo_inputs_t;
        signal fifo_full_140097941553392: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941553392: core_fifo_inputs_t;
        signal outputs_full_140097941553392: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941553448: core_fifo_inputs_t;
        signal fifo_full_140097941553448: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941553448: core_fifo_inputs_t;
        signal outputs_full_140097941553448: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941553504: core_fifo_inputs_t;
        signal fifo_full_140097941553504: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941553504: core_fifo_inputs_t;
        signal outputs_full_140097941553504: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941553560: core_fifo_inputs_t;
        signal fifo_full_140097941553560: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941553560: core_fifo_inputs_t;
        signal outputs_full_140097941553560: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941553616: core_fifo_inputs_t;
        signal fifo_full_140097941553616: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941553616: core_fifo_inputs_t;
        signal outputs_full_140097941553616: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941553672: core_fifo_inputs_t;
        signal fifo_full_140097941553672: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941553672: core_fifo_inputs_t;
        signal outputs_full_140097941553672: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941553728: core_fifo_inputs_t;
        signal fifo_full_140097941553728: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941553728: core_fifo_inputs_t;
        signal outputs_full_140097941553728: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941553784: core_fifo_inputs_t;
        signal fifo_full_140097941553784: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941553784: core_fifo_inputs_t;
        signal outputs_full_140097941553784: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941553840: core_fifo_inputs_t;
        signal fifo_full_140097941553840: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941553840: core_fifo_inputs_t;
        signal outputs_full_140097941553840: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941553896: core_fifo_inputs_t;
        signal fifo_full_140097941553896: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941553896: core_fifo_inputs_t;
        signal outputs_full_140097941553896: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941553952: core_fifo_inputs_t;
        signal fifo_full_140097941553952: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941553952: core_fifo_inputs_t;
        signal outputs_full_140097941553952: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941554008: core_fifo_inputs_t;
        signal fifo_full_140097941554008: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941554008: core_fifo_inputs_t;
        signal outputs_full_140097941554008: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941554064: core_fifo_inputs_t;
        signal fifo_full_140097941554064: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941554064: core_fifo_inputs_t;
        signal outputs_full_140097941554064: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941554120: core_fifo_inputs_t;
        signal fifo_full_140097941554120: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941554120: core_fifo_inputs_t;
        signal outputs_full_140097941554120: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941554176: core_fifo_inputs_t;
        signal fifo_full_140097941554176: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941554176: core_fifo_inputs_t;
        signal outputs_full_140097941554176: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941554232: core_fifo_inputs_t;
        signal fifo_full_140097941554232: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941554232: core_fifo_inputs_t;
        signal outputs_full_140097941554232: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941554288: core_fifo_inputs_t;
        signal fifo_full_140097941554288: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941554288: core_fifo_inputs_t;
        signal outputs_full_140097941554288: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941554344: core_fifo_inputs_t;
        signal fifo_full_140097941554344: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941554344: core_fifo_inputs_t;
        signal outputs_full_140097941554344: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941554400: core_fifo_inputs_t;
        signal fifo_full_140097941554400: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941554400: core_fifo_inputs_t;
        signal outputs_full_140097941554400: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941554456: core_fifo_inputs_t;
        signal fifo_full_140097941554456: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941554456: core_fifo_inputs_t;
        signal outputs_full_140097941554456: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941554512: core_fifo_inputs_t;
        signal fifo_full_140097941554512: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941554512: core_fifo_inputs_t;
        signal outputs_full_140097941554512: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941554568: core_fifo_inputs_t;
        signal fifo_full_140097941554568: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941554568: core_fifo_inputs_t;
        signal outputs_full_140097941554568: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941554624: core_fifo_inputs_t;
        signal fifo_full_140097941554624: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941554624: core_fifo_inputs_t;
        signal outputs_full_140097941554624: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941554680: core_fifo_inputs_t;
        signal fifo_full_140097941554680: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941554680: core_fifo_inputs_t;
        signal outputs_full_140097941554680: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941554736: core_fifo_inputs_t;
        signal fifo_full_140097941554736: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941554736: core_fifo_inputs_t;
        signal outputs_full_140097941554736: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941554792: core_fifo_inputs_t;
        signal fifo_full_140097941554792: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941554792: core_fifo_inputs_t;
        signal outputs_full_140097941554792: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941554848: core_fifo_inputs_t;
        signal fifo_full_140097941554848: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941554848: core_fifo_inputs_t;
        signal outputs_full_140097941554848: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941554904: core_fifo_inputs_t;
        signal fifo_full_140097941554904: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941554904: core_fifo_inputs_t;
        signal outputs_full_140097941554904: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941554960: core_fifo_inputs_t;
        signal fifo_full_140097941554960: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941554960: core_fifo_inputs_t;
        signal outputs_full_140097941554960: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941555016: core_fifo_inputs_t;
        signal fifo_full_140097941555016: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941555016: core_fifo_inputs_t;
        signal outputs_full_140097941555016: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941555072: core_fifo_inputs_t;
        signal fifo_full_140097941555072: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941555072: core_fifo_inputs_t;
        signal outputs_full_140097941555072: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941555128: core_fifo_inputs_t;
        signal fifo_full_140097941555128: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941555128: core_fifo_inputs_t;
        signal outputs_full_140097941555128: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941555184: core_fifo_inputs_t;
        signal fifo_full_140097941555184: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941555184: core_fifo_inputs_t;
        signal outputs_full_140097941555184: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941555240: core_fifo_inputs_t;
        signal fifo_full_140097941555240: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941555240: core_fifo_inputs_t;
        signal outputs_full_140097941555240: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941555296: core_fifo_inputs_t;
        signal fifo_full_140097941555296: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941555296: core_fifo_inputs_t;
        signal outputs_full_140097941555296: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941555352: core_fifo_inputs_t;
        signal fifo_full_140097941555352: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941555352: core_fifo_inputs_t;
        signal outputs_full_140097941555352: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941555408: core_fifo_inputs_t;
        signal fifo_full_140097941555408: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941555408: core_fifo_inputs_t;
        signal outputs_full_140097941555408: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941555464: core_fifo_inputs_t;
        signal fifo_full_140097941555464: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941555464: core_fifo_inputs_t;
        signal outputs_full_140097941555464: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941555520: core_fifo_inputs_t;
        signal fifo_full_140097941555520: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941555520: core_fifo_inputs_t;
        signal outputs_full_140097941555520: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941555576: core_fifo_inputs_t;
        signal fifo_full_140097941555576: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941555576: core_fifo_inputs_t;
        signal outputs_full_140097941555576: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941555632: core_fifo_inputs_t;
        signal fifo_full_140097941555632: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941555632: core_fifo_inputs_t;
        signal outputs_full_140097941555632: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140097941555688: core_fifo_inputs_t;
        signal fifo_full_140097941555688: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140097941555688: core_fifo_inputs_t;
        signal outputs_full_140097941555688: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        

begin

        fifo_inputs_140097944041960 <= fifo_inputs;
        fifo_full <= fifo_full_140097944041960;

        fifo_inputs_140097944041904(0) <= outputs_140097944041960(0);
        outputs_full_140097944041960(0) <= fifo_full_140097944041904(0);
        
        fifo_inputs_140097944042128(0) <= outputs_140097944041904(0);
        outputs_full_140097944041904(0) <= fifo_full_140097944042128(0);
        
        fifo_inputs_140097944042072(0) <= outputs_140097944042128(0);
        outputs_full_140097944042128(0) <= fifo_full_140097944042072(0);
        
        fifo_inputs_140097944042184(0) <= outputs_140097944042072(0);
        outputs_full_140097944042072(0) <= fifo_full_140097944042184(0);
        
        fifo_inputs_140097944042240(0) <= outputs_140097944042184(0);
        outputs_full_140097944042184(0) <= fifo_full_140097944042240(0);
        
        fifo_inputs_140097944042296(0) <= outputs_140097944042240(0);
        outputs_full_140097944042240(0) <= fifo_full_140097944042296(0);
        
        fifo_inputs_140097944042352(0) <= outputs_140097944042296(0);
        outputs_full_140097944042296(0) <= fifo_full_140097944042352(0);
        
        fifo_inputs_140097944042408(0) <= outputs_140097944042352(0);
        outputs_full_140097944042352(0) <= fifo_full_140097944042408(0);
        
        fifo_inputs_140097944042464(0) <= outputs_140097944042408(0);
        outputs_full_140097944042408(0) <= fifo_full_140097944042464(0);
        
        fifo_inputs_140097944042016(0) <= outputs_140097944042464(0);
        outputs_full_140097944042464(0) <= fifo_full_140097944042016(0);
        
        fifo_inputs_140097944042520(0) <= outputs_140097944042016(0);
        outputs_full_140097944042016(0) <= fifo_full_140097944042520(0);
        
        fifo_inputs_140097944042576(0) <= outputs_140097944042520(0);
        outputs_full_140097944042520(0) <= fifo_full_140097944042576(0);
        
        fifo_inputs_140097944042632(0) <= outputs_140097944042576(0);
        outputs_full_140097944042576(0) <= fifo_full_140097944042632(0);
        
        fifo_inputs_140097944042688(0) <= outputs_140097944042632(0);
        outputs_full_140097944042632(0) <= fifo_full_140097944042688(0);
        
        fifo_inputs_140097944042744(0) <= outputs_140097944042688(0);
        outputs_full_140097944042688(0) <= fifo_full_140097944042744(0);
        
        fifo_inputs_140097944042800(0) <= outputs_140097944042744(0);
        outputs_full_140097944042744(0) <= fifo_full_140097944042800(0);
        
        fifo_inputs_140097944042856(0) <= outputs_140097944042800(0);
        outputs_full_140097944042800(0) <= fifo_full_140097944042856(0);
        
        fifo_inputs_140097944042912(0) <= outputs_140097944042856(0);
        outputs_full_140097944042856(0) <= fifo_full_140097944042912(0);
        
        fifo_inputs_140097944042968(0) <= outputs_140097944042912(0);
        outputs_full_140097944042912(0) <= fifo_full_140097944042968(0);
        
        fifo_inputs_140097944043024(0) <= outputs_140097944042968(0);
        outputs_full_140097944042968(0) <= fifo_full_140097944043024(0);
        
        fifo_inputs_140097944043080(0) <= outputs_140097944043024(0);
        outputs_full_140097944043024(0) <= fifo_full_140097944043080(0);
        
        fifo_inputs_140097944043136(0) <= outputs_140097944043080(0);
        outputs_full_140097944043080(0) <= fifo_full_140097944043136(0);
        
        fifo_inputs_140097944043192(0) <= outputs_140097944043136(0);
        outputs_full_140097944043136(0) <= fifo_full_140097944043192(0);
        
        fifo_inputs_140097944043248(0) <= outputs_140097944043192(0);
        outputs_full_140097944043192(0) <= fifo_full_140097944043248(0);
        
        fifo_inputs_140097944043304(0) <= outputs_140097944043248(0);
        outputs_full_140097944043248(0) <= fifo_full_140097944043304(0);
        
        fifo_inputs_140097944043360(0) <= outputs_140097944043304(0);
        outputs_full_140097944043304(0) <= fifo_full_140097944043360(0);
        
        fifo_inputs_140097944043416(0) <= outputs_140097944043360(0);
        outputs_full_140097944043360(0) <= fifo_full_140097944043416(0);
        
        fifo_inputs_140097944043472(0) <= outputs_140097944043416(0);
        outputs_full_140097944043416(0) <= fifo_full_140097944043472(0);
        
        fifo_inputs_140097944076360(0) <= outputs_140097944043472(0);
        outputs_full_140097944043472(0) <= fifo_full_140097944076360(0);
        
        fifo_inputs_140097944076416(0) <= outputs_140097944076360(0);
        outputs_full_140097944076360(0) <= fifo_full_140097944076416(0);
        
        fifo_inputs_140097944076472(0) <= outputs_140097944076416(0);
        outputs_full_140097944076416(0) <= fifo_full_140097944076472(0);
        
        fifo_inputs_140097944076528(0) <= outputs_140097944076472(0);
        outputs_full_140097944076472(0) <= fifo_full_140097944076528(0);
        
        fifo_inputs_140097944076584(0) <= outputs_140097944076528(0);
        outputs_full_140097944076528(0) <= fifo_full_140097944076584(0);
        
        fifo_inputs_140097944076640(0) <= outputs_140097944076584(0);
        outputs_full_140097944076584(0) <= fifo_full_140097944076640(0);
        
        fifo_inputs_140097944076696(0) <= outputs_140097944076640(0);
        outputs_full_140097944076640(0) <= fifo_full_140097944076696(0);
        
        fifo_inputs_140097944076752(0) <= outputs_140097944076696(0);
        outputs_full_140097944076696(0) <= fifo_full_140097944076752(0);
        
        fifo_inputs_140097944076808(0) <= outputs_140097944076752(0);
        outputs_full_140097944076752(0) <= fifo_full_140097944076808(0);
        
        fifo_inputs_140097944076864(0) <= outputs_140097944076808(0);
        outputs_full_140097944076808(0) <= fifo_full_140097944076864(0);
        
        fifo_inputs_140097944076920(0) <= outputs_140097944076864(0);
        outputs_full_140097944076864(0) <= fifo_full_140097944076920(0);
        
        fifo_inputs_140097944076976(0) <= outputs_140097944076920(0);
        outputs_full_140097944076920(0) <= fifo_full_140097944076976(0);
        
        fifo_inputs_140097944077032(0) <= outputs_140097944076976(0);
        outputs_full_140097944076976(0) <= fifo_full_140097944077032(0);
        
        fifo_inputs_140097944077088(0) <= outputs_140097944077032(0);
        outputs_full_140097944077032(0) <= fifo_full_140097944077088(0);
        
        fifo_inputs_140097944077144(0) <= outputs_140097944077088(0);
        outputs_full_140097944077088(0) <= fifo_full_140097944077144(0);
        
        fifo_inputs_140097944077200(0) <= outputs_140097944077144(0);
        outputs_full_140097944077144(0) <= fifo_full_140097944077200(0);
        
        fifo_inputs_140097944077256(0) <= outputs_140097944077200(0);
        outputs_full_140097944077200(0) <= fifo_full_140097944077256(0);
        
        fifo_inputs_140097944077312(0) <= outputs_140097944077256(0);
        outputs_full_140097944077256(0) <= fifo_full_140097944077312(0);
        
        fifo_inputs_140097944077368(0) <= outputs_140097944077312(0);
        outputs_full_140097944077312(0) <= fifo_full_140097944077368(0);
        
        fifo_inputs_140097944077424(0) <= outputs_140097944077368(0);
        outputs_full_140097944077368(0) <= fifo_full_140097944077424(0);
        
        fifo_inputs_140097944077480(0) <= outputs_140097944077424(0);
        outputs_full_140097944077424(0) <= fifo_full_140097944077480(0);
        
        fifo_inputs_140097944077536(0) <= outputs_140097944077480(0);
        outputs_full_140097944077480(0) <= fifo_full_140097944077536(0);
        
        fifo_inputs_140097944077592(0) <= outputs_140097944077536(0);
        outputs_full_140097944077536(0) <= fifo_full_140097944077592(0);
        
        fifo_inputs_140097944077648(0) <= outputs_140097944077592(0);
        outputs_full_140097944077592(0) <= fifo_full_140097944077648(0);
        
        fifo_inputs_140097944077704(0) <= outputs_140097944077648(0);
        outputs_full_140097944077648(0) <= fifo_full_140097944077704(0);
        
        fifo_inputs_140097944077760(0) <= outputs_140097944077704(0);
        outputs_full_140097944077704(0) <= fifo_full_140097944077760(0);
        
        fifo_inputs_140097944077816(0) <= outputs_140097944077760(0);
        outputs_full_140097944077760(0) <= fifo_full_140097944077816(0);
        
        fifo_inputs_140097944077872(0) <= outputs_140097944077816(0);
        outputs_full_140097944077816(0) <= fifo_full_140097944077872(0);
        
        fifo_inputs_140097944077928(0) <= outputs_140097944077872(0);
        outputs_full_140097944077872(0) <= fifo_full_140097944077928(0);
        
        fifo_inputs_140097944077984(0) <= outputs_140097944077928(0);
        outputs_full_140097944077928(0) <= fifo_full_140097944077984(0);
        
        fifo_inputs_140097944078040(0) <= outputs_140097944077984(0);
        outputs_full_140097944077984(0) <= fifo_full_140097944078040(0);
        
        fifo_inputs_140097944078096(0) <= outputs_140097944078040(0);
        outputs_full_140097944078040(0) <= fifo_full_140097944078096(0);
        
        fifo_inputs_140097944078152(0) <= outputs_140097944078096(0);
        outputs_full_140097944078096(0) <= fifo_full_140097944078152(0);
        
        fifo_inputs_140097944078208(0) <= outputs_140097944078152(0);
        outputs_full_140097944078152(0) <= fifo_full_140097944078208(0);
        
        fifo_inputs_140097944078264(0) <= outputs_140097944078208(0);
        outputs_full_140097944078208(0) <= fifo_full_140097944078264(0);
        
        fifo_inputs_140097944078320(0) <= outputs_140097944078264(0);
        outputs_full_140097944078264(0) <= fifo_full_140097944078320(0);
        
        fifo_inputs_140097944078376(0) <= outputs_140097944078320(0);
        outputs_full_140097944078320(0) <= fifo_full_140097944078376(0);
        
        fifo_inputs_140097944078432(0) <= outputs_140097944078376(0);
        outputs_full_140097944078376(0) <= fifo_full_140097944078432(0);
        
        fifo_inputs_140097944078488(0) <= outputs_140097944078432(0);
        outputs_full_140097944078432(0) <= fifo_full_140097944078488(0);
        
        fifo_inputs_140097944078544(0) <= outputs_140097944078488(0);
        outputs_full_140097944078488(0) <= fifo_full_140097944078544(0);
        
        fifo_inputs_140097944078600(0) <= outputs_140097944078544(0);
        outputs_full_140097944078544(0) <= fifo_full_140097944078600(0);
        
        fifo_inputs_140097944078656(0) <= outputs_140097944078600(0);
        outputs_full_140097944078600(0) <= fifo_full_140097944078656(0);
        
        fifo_inputs_140097944078712(0) <= outputs_140097944078656(0);
        outputs_full_140097944078656(0) <= fifo_full_140097944078712(0);
        
        fifo_inputs_140097944078768(0) <= outputs_140097944078712(0);
        outputs_full_140097944078712(0) <= fifo_full_140097944078768(0);
        
        fifo_inputs_140097944078824(0) <= outputs_140097944078768(0);
        outputs_full_140097944078768(0) <= fifo_full_140097944078824(0);
        
        fifo_inputs_140097944078880(0) <= outputs_140097944078824(0);
        outputs_full_140097944078824(0) <= fifo_full_140097944078880(0);
        
        fifo_inputs_140097944078936(0) <= outputs_140097944078880(0);
        outputs_full_140097944078880(0) <= fifo_full_140097944078936(0);
        
        fifo_inputs_140097944078992(0) <= outputs_140097944078936(0);
        outputs_full_140097944078936(0) <= fifo_full_140097944078992(0);
        
        fifo_inputs_140097944079048(0) <= outputs_140097944078992(0);
        outputs_full_140097944078992(0) <= fifo_full_140097944079048(0);
        
        fifo_inputs_140097944079104(0) <= outputs_140097944079048(0);
        outputs_full_140097944079048(0) <= fifo_full_140097944079104(0);
        
        fifo_inputs_140097944079160(0) <= outputs_140097944079104(0);
        outputs_full_140097944079104(0) <= fifo_full_140097944079160(0);
        
        fifo_inputs_140097944079216(0) <= outputs_140097944079160(0);
        outputs_full_140097944079160(0) <= fifo_full_140097944079216(0);
        
        fifo_inputs_140097944079272(0) <= outputs_140097944079216(0);
        outputs_full_140097944079216(0) <= fifo_full_140097944079272(0);
        
        fifo_inputs_140097944079328(0) <= outputs_140097944079272(0);
        outputs_full_140097944079272(0) <= fifo_full_140097944079328(0);
        
        fifo_inputs_140097944079384(0) <= outputs_140097944079328(0);
        outputs_full_140097944079328(0) <= fifo_full_140097944079384(0);
        
        fifo_inputs_140097944079440(0) <= outputs_140097944079384(0);
        outputs_full_140097944079384(0) <= fifo_full_140097944079440(0);
        
        fifo_inputs_140097944079496(0) <= outputs_140097944079440(0);
        outputs_full_140097944079440(0) <= fifo_full_140097944079496(0);
        
        fifo_inputs_140097944079552(0) <= outputs_140097944079496(0);
        outputs_full_140097944079496(0) <= fifo_full_140097944079552(0);
        
        fifo_inputs_140097944079608(0) <= outputs_140097944079552(0);
        outputs_full_140097944079552(0) <= fifo_full_140097944079608(0);
        
        fifo_inputs_140097944079664(0) <= outputs_140097944079608(0);
        outputs_full_140097944079608(0) <= fifo_full_140097944079664(0);
        
        fifo_inputs_140097944079720(0) <= outputs_140097944079664(0);
        outputs_full_140097944079664(0) <= fifo_full_140097944079720(0);
        
        fifo_inputs_140097944079776(0) <= outputs_140097944079720(0);
        outputs_full_140097944079720(0) <= fifo_full_140097944079776(0);
        
        fifo_inputs_140097944079832(0) <= outputs_140097944079776(0);
        outputs_full_140097944079776(0) <= fifo_full_140097944079832(0);
        
        fifo_inputs_140097944079888(0) <= outputs_140097944079832(0);
        outputs_full_140097944079832(0) <= fifo_full_140097944079888(0);
        
        fifo_inputs_140097944079944(0) <= outputs_140097944079888(0);
        outputs_full_140097944079888(0) <= fifo_full_140097944079944(0);
        
        fifo_inputs_140097944080000(0) <= outputs_140097944079944(0);
        outputs_full_140097944079944(0) <= fifo_full_140097944080000(0);
        
        fifo_inputs_140097944080056(0) <= outputs_140097944080000(0);
        outputs_full_140097944080000(0) <= fifo_full_140097944080056(0);
        
        fifo_inputs_140097944080112(0) <= outputs_140097944080056(0);
        outputs_full_140097944080056(0) <= fifo_full_140097944080112(0);
        
        fifo_inputs_140097944080168(0) <= outputs_140097944080112(0);
        outputs_full_140097944080112(0) <= fifo_full_140097944080168(0);
        
        fifo_inputs_140097944080224(0) <= outputs_140097944080168(0);
        outputs_full_140097944080168(0) <= fifo_full_140097944080224(0);
        
        fifo_inputs_140097944080280(0) <= outputs_140097944080224(0);
        outputs_full_140097944080224(0) <= fifo_full_140097944080280(0);
        
        fifo_inputs_140097944080336(0) <= outputs_140097944080280(0);
        outputs_full_140097944080280(0) <= fifo_full_140097944080336(0);
        
        fifo_inputs_140097944096840(0) <= outputs_140097944080336(0);
        outputs_full_140097944080336(0) <= fifo_full_140097944096840(0);
        
        fifo_inputs_140097944096896(0) <= outputs_140097944096840(0);
        outputs_full_140097944096840(0) <= fifo_full_140097944096896(0);
        
        fifo_inputs_140097944096952(0) <= outputs_140097944096896(0);
        outputs_full_140097944096896(0) <= fifo_full_140097944096952(0);
        
        fifo_inputs_140097944097008(0) <= outputs_140097944096952(0);
        outputs_full_140097944096952(0) <= fifo_full_140097944097008(0);
        
        fifo_inputs_140097944097064(0) <= outputs_140097944097008(0);
        outputs_full_140097944097008(0) <= fifo_full_140097944097064(0);
        
        fifo_inputs_140097944097120(0) <= outputs_140097944097064(0);
        outputs_full_140097944097064(0) <= fifo_full_140097944097120(0);
        
        fifo_inputs_140097944097176(0) <= outputs_140097944097120(0);
        outputs_full_140097944097120(0) <= fifo_full_140097944097176(0);
        
        fifo_inputs_140097944097232(0) <= outputs_140097944097176(0);
        outputs_full_140097944097176(0) <= fifo_full_140097944097232(0);
        
        fifo_inputs_140097944097288(0) <= outputs_140097944097232(0);
        outputs_full_140097944097232(0) <= fifo_full_140097944097288(0);
        
        fifo_inputs_140097944097344(0) <= outputs_140097944097288(0);
        outputs_full_140097944097288(0) <= fifo_full_140097944097344(0);
        
        fifo_inputs_140097944097400(0) <= outputs_140097944097344(0);
        outputs_full_140097944097344(0) <= fifo_full_140097944097400(0);
        
        fifo_inputs_140097944097456(0) <= outputs_140097944097400(0);
        outputs_full_140097944097400(0) <= fifo_full_140097944097456(0);
        
        fifo_inputs_140097944097512(0) <= outputs_140097944097456(0);
        outputs_full_140097944097456(0) <= fifo_full_140097944097512(0);
        
        fifo_inputs_140097944097568(0) <= outputs_140097944097512(0);
        outputs_full_140097944097512(0) <= fifo_full_140097944097568(0);
        
        fifo_inputs_140097944097624(0) <= outputs_140097944097568(0);
        outputs_full_140097944097568(0) <= fifo_full_140097944097624(0);
        
        fifo_inputs_140097944097680(0) <= outputs_140097944097624(0);
        outputs_full_140097944097624(0) <= fifo_full_140097944097680(0);
        
        fifo_inputs_140097944097736(0) <= outputs_140097944097680(0);
        outputs_full_140097944097680(0) <= fifo_full_140097944097736(0);
        
        fifo_inputs_140097944097792(0) <= outputs_140097944097736(0);
        outputs_full_140097944097736(0) <= fifo_full_140097944097792(0);
        
        fifo_inputs_140097944097848(0) <= outputs_140097944097792(0);
        outputs_full_140097944097792(0) <= fifo_full_140097944097848(0);
        
        fifo_inputs_140097944097904(0) <= outputs_140097944097848(0);
        outputs_full_140097944097848(0) <= fifo_full_140097944097904(0);
        
        fifo_inputs_140097944097960(0) <= outputs_140097944097904(0);
        outputs_full_140097944097904(0) <= fifo_full_140097944097960(0);
        
        fifo_inputs_140097944098016(0) <= outputs_140097944097960(0);
        outputs_full_140097944097960(0) <= fifo_full_140097944098016(0);
        
        fifo_inputs_140097944098072(0) <= outputs_140097944098016(0);
        outputs_full_140097944098016(0) <= fifo_full_140097944098072(0);
        
        fifo_inputs_140097944098128(0) <= outputs_140097944098072(0);
        outputs_full_140097944098072(0) <= fifo_full_140097944098128(0);
        
        fifo_inputs_140097944098184(0) <= outputs_140097944098128(0);
        outputs_full_140097944098128(0) <= fifo_full_140097944098184(0);
        
        fifo_inputs_140097944098240(0) <= outputs_140097944098184(0);
        outputs_full_140097944098184(0) <= fifo_full_140097944098240(0);
        
        fifo_inputs_140097944098296(0) <= outputs_140097944098240(0);
        outputs_full_140097944098240(0) <= fifo_full_140097944098296(0);
        
        fifo_inputs_140097944098352(0) <= outputs_140097944098296(0);
        outputs_full_140097944098296(0) <= fifo_full_140097944098352(0);
        
        fifo_inputs_140097944098408(0) <= outputs_140097944098352(0);
        outputs_full_140097944098352(0) <= fifo_full_140097944098408(0);
        
        fifo_inputs_140097944098464(0) <= outputs_140097944098408(0);
        outputs_full_140097944098408(0) <= fifo_full_140097944098464(0);
        
        fifo_inputs_140097944098520(0) <= outputs_140097944098464(0);
        outputs_full_140097944098464(0) <= fifo_full_140097944098520(0);
        
        fifo_inputs_140097944098576(0) <= outputs_140097944098520(0);
        outputs_full_140097944098520(0) <= fifo_full_140097944098576(0);
        
        fifo_inputs_140097944098632(0) <= outputs_140097944098576(0);
        outputs_full_140097944098576(0) <= fifo_full_140097944098632(0);
        
        fifo_inputs_140097944098688(0) <= outputs_140097944098632(0);
        outputs_full_140097944098632(0) <= fifo_full_140097944098688(0);
        
        fifo_inputs_140097944098744(0) <= outputs_140097944098688(0);
        outputs_full_140097944098688(0) <= fifo_full_140097944098744(0);
        
        fifo_inputs_140097944098800(0) <= outputs_140097944098744(0);
        outputs_full_140097944098744(0) <= fifo_full_140097944098800(0);
        
        fifo_inputs_140097944098856(0) <= outputs_140097944098800(0);
        outputs_full_140097944098800(0) <= fifo_full_140097944098856(0);
        
        fifo_inputs_140097944098912(0) <= outputs_140097944098856(0);
        outputs_full_140097944098856(0) <= fifo_full_140097944098912(0);
        
        fifo_inputs_140097944098968(0) <= outputs_140097944098912(0);
        outputs_full_140097944098912(0) <= fifo_full_140097944098968(0);
        
        fifo_inputs_140097944099024(0) <= outputs_140097944098968(0);
        outputs_full_140097944098968(0) <= fifo_full_140097944099024(0);
        
        fifo_inputs_140097944099080(0) <= outputs_140097944099024(0);
        outputs_full_140097944099024(0) <= fifo_full_140097944099080(0);
        
        fifo_inputs_140097944099136(0) <= outputs_140097944099080(0);
        outputs_full_140097944099080(0) <= fifo_full_140097944099136(0);
        
        fifo_inputs_140097944099192(0) <= outputs_140097944099136(0);
        outputs_full_140097944099136(0) <= fifo_full_140097944099192(0);
        
        fifo_inputs_140097944099248(0) <= outputs_140097944099192(0);
        outputs_full_140097944099192(0) <= fifo_full_140097944099248(0);
        
        fifo_inputs_140097944099304(0) <= outputs_140097944099248(0);
        outputs_full_140097944099248(0) <= fifo_full_140097944099304(0);
        
        fifo_inputs_140097944099360(0) <= outputs_140097944099304(0);
        outputs_full_140097944099304(0) <= fifo_full_140097944099360(0);
        
        fifo_inputs_140097944099416(0) <= outputs_140097944099360(0);
        outputs_full_140097944099360(0) <= fifo_full_140097944099416(0);
        
        fifo_inputs_140097944099472(0) <= outputs_140097944099416(0);
        outputs_full_140097944099416(0) <= fifo_full_140097944099472(0);
        
        fifo_inputs_140097944099528(0) <= outputs_140097944099472(0);
        outputs_full_140097944099472(0) <= fifo_full_140097944099528(0);
        
        fifo_inputs_140097965543496(0) <= outputs_140097944099528(0);
        outputs_full_140097944099528(0) <= fifo_full_140097965543496(0);
        
        fifo_inputs_140097944041736(0) <= outputs_140097965543496(0);
        outputs_full_140097965543496(0) <= fifo_full_140097944041736(0);
        
        fifo_inputs_140097944041624(0) <= outputs_140097944041736(0);
        outputs_full_140097944041736(0) <= fifo_full_140097944041624(0);
        
        fifo_inputs_140097944041568(0) <= outputs_140097944041624(0);
        outputs_full_140097944041624(0) <= fifo_full_140097944041568(0);
        
        fifo_inputs_140097944041792(0) <= outputs_140097944041568(0);
        outputs_full_140097944041568(0) <= fifo_full_140097944041792(0);
        
        fifo_inputs_140097944041456(0) <= outputs_140097944041792(0);
        outputs_full_140097944041792(0) <= fifo_full_140097944041456(0);
        
        fifo_inputs_140097944099584(0) <= outputs_140097944041456(0);
        outputs_full_140097944041456(0) <= fifo_full_140097944099584(0);
        
        fifo_inputs_140097944099640(0) <= outputs_140097944099584(0);
        outputs_full_140097944099584(0) <= fifo_full_140097944099640(0);
        
        fifo_inputs_140097944099696(0) <= outputs_140097944099640(0);
        outputs_full_140097944099640(0) <= fifo_full_140097944099696(0);
        
        fifo_inputs_140097944099752(0) <= outputs_140097944099696(0);
        outputs_full_140097944099696(0) <= fifo_full_140097944099752(0);
        
        fifo_inputs_140097944099808(0) <= outputs_140097944099752(0);
        outputs_full_140097944099752(0) <= fifo_full_140097944099808(0);
        
        fifo_inputs_140097944099864(0) <= outputs_140097944099808(0);
        outputs_full_140097944099808(0) <= fifo_full_140097944099864(0);
        
        fifo_inputs_140097944099920(0) <= outputs_140097944099864(0);
        outputs_full_140097944099864(0) <= fifo_full_140097944099920(0);
        
        fifo_inputs_140097944099976(0) <= outputs_140097944099920(0);
        outputs_full_140097944099920(0) <= fifo_full_140097944099976(0);
        
        fifo_inputs_140097944100032(0) <= outputs_140097944099976(0);
        outputs_full_140097944099976(0) <= fifo_full_140097944100032(0);
        
        fifo_inputs_140097944100088(0) <= outputs_140097944100032(0);
        outputs_full_140097944100032(0) <= fifo_full_140097944100088(0);
        
        fifo_inputs_140097944100144(0) <= outputs_140097944100088(0);
        outputs_full_140097944100088(0) <= fifo_full_140097944100144(0);
        
        fifo_inputs_140097944100200(0) <= outputs_140097944100144(0);
        outputs_full_140097944100144(0) <= fifo_full_140097944100200(0);
        
        fifo_inputs_140097944100256(0) <= outputs_140097944100200(0);
        outputs_full_140097944100200(0) <= fifo_full_140097944100256(0);
        
        fifo_inputs_140097944100312(0) <= outputs_140097944100256(0);
        outputs_full_140097944100256(0) <= fifo_full_140097944100312(0);
        
        fifo_inputs_140097944100368(0) <= outputs_140097944100312(0);
        outputs_full_140097944100312(0) <= fifo_full_140097944100368(0);
        
        fifo_inputs_140097944100424(0) <= outputs_140097944100368(0);
        outputs_full_140097944100368(0) <= fifo_full_140097944100424(0);
        
        fifo_inputs_140097944100480(0) <= outputs_140097944100424(0);
        outputs_full_140097944100424(0) <= fifo_full_140097944100480(0);
        
        fifo_inputs_140097944100536(0) <= outputs_140097944100480(0);
        outputs_full_140097944100480(0) <= fifo_full_140097944100536(0);
        
        fifo_inputs_140097944100592(0) <= outputs_140097944100536(0);
        outputs_full_140097944100536(0) <= fifo_full_140097944100592(0);
        
        fifo_inputs_140097944100648(0) <= outputs_140097944100592(0);
        outputs_full_140097944100592(0) <= fifo_full_140097944100648(0);
        
        fifo_inputs_140097944100704(0) <= outputs_140097944100648(0);
        outputs_full_140097944100648(0) <= fifo_full_140097944100704(0);
        
        fifo_inputs_140097944100760(0) <= outputs_140097944100704(0);
        outputs_full_140097944100704(0) <= fifo_full_140097944100760(0);
        
        fifo_inputs_140097944100816(0) <= outputs_140097944100760(0);
        outputs_full_140097944100760(0) <= fifo_full_140097944100816(0);
        
        fifo_inputs_140097944113224(0) <= outputs_140097944100816(0);
        outputs_full_140097944100816(0) <= fifo_full_140097944113224(0);
        
        fifo_inputs_140097944113280(0) <= outputs_140097944113224(0);
        outputs_full_140097944113224(0) <= fifo_full_140097944113280(0);
        
        fifo_inputs_140097944113336(0) <= outputs_140097944113280(0);
        outputs_full_140097944113280(0) <= fifo_full_140097944113336(0);
        
        fifo_inputs_140097944113392(0) <= outputs_140097944113336(0);
        outputs_full_140097944113336(0) <= fifo_full_140097944113392(0);
        
        fifo_inputs_140097944113448(0) <= outputs_140097944113392(0);
        outputs_full_140097944113392(0) <= fifo_full_140097944113448(0);
        
        fifo_inputs_140097944113504(0) <= outputs_140097944113448(0);
        outputs_full_140097944113448(0) <= fifo_full_140097944113504(0);
        
        fifo_inputs_140097944113560(0) <= outputs_140097944113504(0);
        outputs_full_140097944113504(0) <= fifo_full_140097944113560(0);
        
        fifo_inputs_140097944113616(0) <= outputs_140097944113560(0);
        outputs_full_140097944113560(0) <= fifo_full_140097944113616(0);
        
        fifo_inputs_140097944113672(0) <= outputs_140097944113616(0);
        outputs_full_140097944113616(0) <= fifo_full_140097944113672(0);
        
        fifo_inputs_140097944113728(0) <= outputs_140097944113672(0);
        outputs_full_140097944113672(0) <= fifo_full_140097944113728(0);
        
        fifo_inputs_140097944113784(0) <= outputs_140097944113728(0);
        outputs_full_140097944113728(0) <= fifo_full_140097944113784(0);
        
        fifo_inputs_140097944113840(0) <= outputs_140097944113784(0);
        outputs_full_140097944113784(0) <= fifo_full_140097944113840(0);
        
        fifo_inputs_140097944113896(0) <= outputs_140097944113840(0);
        outputs_full_140097944113840(0) <= fifo_full_140097944113896(0);
        
        fifo_inputs_140097944113952(0) <= outputs_140097944113896(0);
        outputs_full_140097944113896(0) <= fifo_full_140097944113952(0);
        
        fifo_inputs_140097944114008(0) <= outputs_140097944113952(0);
        outputs_full_140097944113952(0) <= fifo_full_140097944114008(0);
        
        fifo_inputs_140097944114064(0) <= outputs_140097944114008(0);
        outputs_full_140097944114008(0) <= fifo_full_140097944114064(0);
        
        fifo_inputs_140097944114120(0) <= outputs_140097944114064(0);
        outputs_full_140097944114064(0) <= fifo_full_140097944114120(0);
        
        fifo_inputs_140097944114176(0) <= outputs_140097944114120(0);
        outputs_full_140097944114120(0) <= fifo_full_140097944114176(0);
        
        fifo_inputs_140097944114232(0) <= outputs_140097944114176(0);
        outputs_full_140097944114176(0) <= fifo_full_140097944114232(0);
        
        fifo_inputs_140097944114288(0) <= outputs_140097944114232(0);
        outputs_full_140097944114232(0) <= fifo_full_140097944114288(0);
        
        fifo_inputs_140097944114344(0) <= outputs_140097944114288(0);
        outputs_full_140097944114288(0) <= fifo_full_140097944114344(0);
        
        fifo_inputs_140097944114400(0) <= outputs_140097944114344(0);
        outputs_full_140097944114344(0) <= fifo_full_140097944114400(0);
        
        fifo_inputs_140097944114456(0) <= outputs_140097944114400(0);
        outputs_full_140097944114400(0) <= fifo_full_140097944114456(0);
        
        fifo_inputs_140097944114512(0) <= outputs_140097944114456(0);
        outputs_full_140097944114456(0) <= fifo_full_140097944114512(0);
        
        fifo_inputs_140097944114568(0) <= outputs_140097944114512(0);
        outputs_full_140097944114512(0) <= fifo_full_140097944114568(0);
        
        fifo_inputs_140097944114624(0) <= outputs_140097944114568(0);
        outputs_full_140097944114568(0) <= fifo_full_140097944114624(0);
        
        fifo_inputs_140097944114680(0) <= outputs_140097944114624(0);
        outputs_full_140097944114624(0) <= fifo_full_140097944114680(0);
        
        fifo_inputs_140097944114736(0) <= outputs_140097944114680(0);
        outputs_full_140097944114680(0) <= fifo_full_140097944114736(0);
        
        fifo_inputs_140097944114792(0) <= outputs_140097944114736(0);
        outputs_full_140097944114736(0) <= fifo_full_140097944114792(0);
        
        fifo_inputs_140097944114848(0) <= outputs_140097944114792(0);
        outputs_full_140097944114792(0) <= fifo_full_140097944114848(0);
        
        fifo_inputs_140097944114904(0) <= outputs_140097944114848(0);
        outputs_full_140097944114848(0) <= fifo_full_140097944114904(0);
        
        fifo_inputs_140097944114960(0) <= outputs_140097944114904(0);
        outputs_full_140097944114904(0) <= fifo_full_140097944114960(0);
        
        fifo_inputs_140097944115016(0) <= outputs_140097944114960(0);
        outputs_full_140097944114960(0) <= fifo_full_140097944115016(0);
        
        fifo_inputs_140097944115072(0) <= outputs_140097944115016(0);
        outputs_full_140097944115016(0) <= fifo_full_140097944115072(0);
        
        fifo_inputs_140097944115128(0) <= outputs_140097944115072(0);
        outputs_full_140097944115072(0) <= fifo_full_140097944115128(0);
        
        fifo_inputs_140097944115184(0) <= outputs_140097944115128(0);
        outputs_full_140097944115128(0) <= fifo_full_140097944115184(0);
        
        fifo_inputs_140097944115240(0) <= outputs_140097944115184(0);
        outputs_full_140097944115184(0) <= fifo_full_140097944115240(0);
        
        fifo_inputs_140097944115296(0) <= outputs_140097944115240(0);
        outputs_full_140097944115240(0) <= fifo_full_140097944115296(0);
        
        fifo_inputs_140097944115352(0) <= outputs_140097944115296(0);
        outputs_full_140097944115296(0) <= fifo_full_140097944115352(0);
        
        fifo_inputs_140097944115408(0) <= outputs_140097944115352(0);
        outputs_full_140097944115352(0) <= fifo_full_140097944115408(0);
        
        fifo_inputs_140097944115464(0) <= outputs_140097944115408(0);
        outputs_full_140097944115408(0) <= fifo_full_140097944115464(0);
        
        fifo_inputs_140097944115520(0) <= outputs_140097944115464(0);
        outputs_full_140097944115464(0) <= fifo_full_140097944115520(0);
        
        fifo_inputs_140097944115576(0) <= outputs_140097944115520(0);
        outputs_full_140097944115520(0) <= fifo_full_140097944115576(0);
        
        fifo_inputs_140097944115632(0) <= outputs_140097944115576(0);
        outputs_full_140097944115576(0) <= fifo_full_140097944115632(0);
        
        fifo_inputs_140097944115688(0) <= outputs_140097944115632(0);
        outputs_full_140097944115632(0) <= fifo_full_140097944115688(0);
        
        fifo_inputs_140097944115744(0) <= outputs_140097944115688(0);
        outputs_full_140097944115688(0) <= fifo_full_140097944115744(0);
        
        fifo_inputs_140097944115800(0) <= outputs_140097944115744(0);
        outputs_full_140097944115744(0) <= fifo_full_140097944115800(0);
        
        fifo_inputs_140097944115856(0) <= outputs_140097944115800(0);
        outputs_full_140097944115800(0) <= fifo_full_140097944115856(0);
        
        fifo_inputs_140097944115912(0) <= outputs_140097944115856(0);
        outputs_full_140097944115856(0) <= fifo_full_140097944115912(0);
        
        fifo_inputs_140097944115968(0) <= outputs_140097944115912(0);
        outputs_full_140097944115912(0) <= fifo_full_140097944115968(0);
        
        fifo_inputs_140097944116024(0) <= outputs_140097944115968(0);
        outputs_full_140097944115968(0) <= fifo_full_140097944116024(0);
        
        fifo_inputs_140097944116080(0) <= outputs_140097944116024(0);
        outputs_full_140097944116024(0) <= fifo_full_140097944116080(0);
        
        fifo_inputs_140097944116136(0) <= outputs_140097944116080(0);
        outputs_full_140097944116080(0) <= fifo_full_140097944116136(0);
        
        fifo_inputs_140097944116192(0) <= outputs_140097944116136(0);
        outputs_full_140097944116136(0) <= fifo_full_140097944116192(0);
        
        fifo_inputs_140097944116248(0) <= outputs_140097944116192(0);
        outputs_full_140097944116192(0) <= fifo_full_140097944116248(0);
        
        fifo_inputs_140097944116304(0) <= outputs_140097944116248(0);
        outputs_full_140097944116248(0) <= fifo_full_140097944116304(0);
        
        fifo_inputs_140097944116360(0) <= outputs_140097944116304(0);
        outputs_full_140097944116304(0) <= fifo_full_140097944116360(0);
        
        fifo_inputs_140097944116416(0) <= outputs_140097944116360(0);
        outputs_full_140097944116360(0) <= fifo_full_140097944116416(0);
        
        fifo_inputs_140097944116472(0) <= outputs_140097944116416(0);
        outputs_full_140097944116416(0) <= fifo_full_140097944116472(0);
        
        fifo_inputs_140097944116528(0) <= outputs_140097944116472(0);
        outputs_full_140097944116472(0) <= fifo_full_140097944116528(0);
        
        fifo_inputs_140097944116584(0) <= outputs_140097944116528(0);
        outputs_full_140097944116528(0) <= fifo_full_140097944116584(0);
        
        fifo_inputs_140097944116640(0) <= outputs_140097944116584(0);
        outputs_full_140097944116584(0) <= fifo_full_140097944116640(0);
        
        fifo_inputs_140097944116696(0) <= outputs_140097944116640(0);
        outputs_full_140097944116640(0) <= fifo_full_140097944116696(0);
        
        fifo_inputs_140097944116752(0) <= outputs_140097944116696(0);
        outputs_full_140097944116696(0) <= fifo_full_140097944116752(0);
        
        fifo_inputs_140097944116808(0) <= outputs_140097944116752(0);
        outputs_full_140097944116752(0) <= fifo_full_140097944116808(0);
        
        fifo_inputs_140097944116864(0) <= outputs_140097944116808(0);
        outputs_full_140097944116808(0) <= fifo_full_140097944116864(0);
        
        fifo_inputs_140097944116920(0) <= outputs_140097944116864(0);
        outputs_full_140097944116864(0) <= fifo_full_140097944116920(0);
        
        fifo_inputs_140097944116976(0) <= outputs_140097944116920(0);
        outputs_full_140097944116920(0) <= fifo_full_140097944116976(0);
        
        fifo_inputs_140097944117032(0) <= outputs_140097944116976(0);
        outputs_full_140097944116976(0) <= fifo_full_140097944117032(0);
        
        fifo_inputs_140097944117088(0) <= outputs_140097944117032(0);
        outputs_full_140097944117032(0) <= fifo_full_140097944117088(0);
        
        fifo_inputs_140097944117144(0) <= outputs_140097944117088(0);
        outputs_full_140097944117088(0) <= fifo_full_140097944117144(0);
        
        fifo_inputs_140097944117200(0) <= outputs_140097944117144(0);
        outputs_full_140097944117144(0) <= fifo_full_140097944117200(0);
        
        fifo_inputs_140097944125512(0) <= outputs_140097944117200(0);
        outputs_full_140097944117200(0) <= fifo_full_140097944125512(0);
        
        fifo_inputs_140097944125568(0) <= outputs_140097944125512(0);
        outputs_full_140097944125512(0) <= fifo_full_140097944125568(0);
        
        fifo_inputs_140097944125624(0) <= outputs_140097944125568(0);
        outputs_full_140097944125568(0) <= fifo_full_140097944125624(0);
        
        fifo_inputs_140097944125680(0) <= outputs_140097944125624(0);
        outputs_full_140097944125624(0) <= fifo_full_140097944125680(0);
        
        fifo_inputs_140097944125736(0) <= outputs_140097944125680(0);
        outputs_full_140097944125680(0) <= fifo_full_140097944125736(0);
        
        fifo_inputs_140097944125792(0) <= outputs_140097944125736(0);
        outputs_full_140097944125736(0) <= fifo_full_140097944125792(0);
        
        fifo_inputs_140097944125848(0) <= outputs_140097944125792(0);
        outputs_full_140097944125792(0) <= fifo_full_140097944125848(0);
        
        fifo_inputs_140097944125904(0) <= outputs_140097944125848(0);
        outputs_full_140097944125848(0) <= fifo_full_140097944125904(0);
        
        fifo_inputs_140097944125960(0) <= outputs_140097944125904(0);
        outputs_full_140097944125904(0) <= fifo_full_140097944125960(0);
        
        fifo_inputs_140097944126016(0) <= outputs_140097944125960(0);
        outputs_full_140097944125960(0) <= fifo_full_140097944126016(0);
        
        fifo_inputs_140097944126072(0) <= outputs_140097944126016(0);
        outputs_full_140097944126016(0) <= fifo_full_140097944126072(0);
        
        fifo_inputs_140097944126128(0) <= outputs_140097944126072(0);
        outputs_full_140097944126072(0) <= fifo_full_140097944126128(0);
        
        fifo_inputs_140097944126184(0) <= outputs_140097944126128(0);
        outputs_full_140097944126128(0) <= fifo_full_140097944126184(0);
        
        fifo_inputs_140097944126240(0) <= outputs_140097944126184(0);
        outputs_full_140097944126184(0) <= fifo_full_140097944126240(0);
        
        fifo_inputs_140097944126296(0) <= outputs_140097944126240(0);
        outputs_full_140097944126240(0) <= fifo_full_140097944126296(0);
        
        fifo_inputs_140097944126352(0) <= outputs_140097944126296(0);
        outputs_full_140097944126296(0) <= fifo_full_140097944126352(0);
        
        fifo_inputs_140097944126408(0) <= outputs_140097944126352(0);
        outputs_full_140097944126352(0) <= fifo_full_140097944126408(0);
        
        fifo_inputs_140097944126464(0) <= outputs_140097944126408(0);
        outputs_full_140097944126408(0) <= fifo_full_140097944126464(0);
        
        fifo_inputs_140097944126520(0) <= outputs_140097944126464(0);
        outputs_full_140097944126464(0) <= fifo_full_140097944126520(0);
        
        fifo_inputs_140097944126576(0) <= outputs_140097944126520(0);
        outputs_full_140097944126520(0) <= fifo_full_140097944126576(0);
        
        fifo_inputs_140097944126632(0) <= outputs_140097944126576(0);
        outputs_full_140097944126576(0) <= fifo_full_140097944126632(0);
        
        fifo_inputs_140097944126688(0) <= outputs_140097944126632(0);
        outputs_full_140097944126632(0) <= fifo_full_140097944126688(0);
        
        fifo_inputs_140097944126744(0) <= outputs_140097944126688(0);
        outputs_full_140097944126688(0) <= fifo_full_140097944126744(0);
        
        fifo_inputs_140097944126800(0) <= outputs_140097944126744(0);
        outputs_full_140097944126744(0) <= fifo_full_140097944126800(0);
        
        fifo_inputs_140097944126856(0) <= outputs_140097944126800(0);
        outputs_full_140097944126800(0) <= fifo_full_140097944126856(0);
        
        fifo_inputs_140097944126912(0) <= outputs_140097944126856(0);
        outputs_full_140097944126856(0) <= fifo_full_140097944126912(0);
        
        fifo_inputs_140097944126968(0) <= outputs_140097944126912(0);
        outputs_full_140097944126912(0) <= fifo_full_140097944126968(0);
        
        fifo_inputs_140097944127024(0) <= outputs_140097944126968(0);
        outputs_full_140097944126968(0) <= fifo_full_140097944127024(0);
        
        fifo_inputs_140097944127080(0) <= outputs_140097944127024(0);
        outputs_full_140097944127024(0) <= fifo_full_140097944127080(0);
        
        fifo_inputs_140097944127136(0) <= outputs_140097944127080(0);
        outputs_full_140097944127080(0) <= fifo_full_140097944127136(0);
        
        fifo_inputs_140097944127192(0) <= outputs_140097944127136(0);
        outputs_full_140097944127136(0) <= fifo_full_140097944127192(0);
        
        fifo_inputs_140097944127248(0) <= outputs_140097944127192(0);
        outputs_full_140097944127192(0) <= fifo_full_140097944127248(0);
        
        fifo_inputs_140097944127304(0) <= outputs_140097944127248(0);
        outputs_full_140097944127248(0) <= fifo_full_140097944127304(0);
        
        fifo_inputs_140097944127360(0) <= outputs_140097944127304(0);
        outputs_full_140097944127304(0) <= fifo_full_140097944127360(0);
        
        fifo_inputs_140097944127416(0) <= outputs_140097944127360(0);
        outputs_full_140097944127360(0) <= fifo_full_140097944127416(0);
        
        fifo_inputs_140097944127472(0) <= outputs_140097944127416(0);
        outputs_full_140097944127416(0) <= fifo_full_140097944127472(0);
        
        fifo_inputs_140097944127528(0) <= outputs_140097944127472(0);
        outputs_full_140097944127472(0) <= fifo_full_140097944127528(0);
        
        fifo_inputs_140097944127584(0) <= outputs_140097944127528(0);
        outputs_full_140097944127528(0) <= fifo_full_140097944127584(0);
        
        fifo_inputs_140097944127640(0) <= outputs_140097944127584(0);
        outputs_full_140097944127584(0) <= fifo_full_140097944127640(0);
        
        fifo_inputs_140097944127696(0) <= outputs_140097944127640(0);
        outputs_full_140097944127640(0) <= fifo_full_140097944127696(0);
        
        fifo_inputs_140097944127752(0) <= outputs_140097944127696(0);
        outputs_full_140097944127696(0) <= fifo_full_140097944127752(0);
        
        fifo_inputs_140097944127808(0) <= outputs_140097944127752(0);
        outputs_full_140097944127752(0) <= fifo_full_140097944127808(0);
        
        fifo_inputs_140097944127864(0) <= outputs_140097944127808(0);
        outputs_full_140097944127808(0) <= fifo_full_140097944127864(0);
        
        fifo_inputs_140097944127920(0) <= outputs_140097944127864(0);
        outputs_full_140097944127864(0) <= fifo_full_140097944127920(0);
        
        fifo_inputs_140097944127976(0) <= outputs_140097944127920(0);
        outputs_full_140097944127920(0) <= fifo_full_140097944127976(0);
        
        fifo_inputs_140097944128032(0) <= outputs_140097944127976(0);
        outputs_full_140097944127976(0) <= fifo_full_140097944128032(0);
        
        fifo_inputs_140097944128088(0) <= outputs_140097944128032(0);
        outputs_full_140097944128032(0) <= fifo_full_140097944128088(0);
        
        fifo_inputs_140097944128144(0) <= outputs_140097944128088(0);
        outputs_full_140097944128088(0) <= fifo_full_140097944128144(0);
        
        fifo_inputs_140097944128200(0) <= outputs_140097944128144(0);
        outputs_full_140097944128144(0) <= fifo_full_140097944128200(0);
        
        fifo_inputs_140097944128256(0) <= outputs_140097944128200(0);
        outputs_full_140097944128200(0) <= fifo_full_140097944128256(0);
        
        fifo_inputs_140097944128312(0) <= outputs_140097944128256(0);
        outputs_full_140097944128256(0) <= fifo_full_140097944128312(0);
        
        fifo_inputs_140097944128368(0) <= outputs_140097944128312(0);
        outputs_full_140097944128312(0) <= fifo_full_140097944128368(0);
        
        fifo_inputs_140097944128424(0) <= outputs_140097944128368(0);
        outputs_full_140097944128368(0) <= fifo_full_140097944128424(0);
        
        fifo_inputs_140097944128480(0) <= outputs_140097944128424(0);
        outputs_full_140097944128424(0) <= fifo_full_140097944128480(0);
        
        fifo_inputs_140097944128536(0) <= outputs_140097944128480(0);
        outputs_full_140097944128480(0) <= fifo_full_140097944128536(0);
        
        fifo_inputs_140097944128592(0) <= outputs_140097944128536(0);
        outputs_full_140097944128536(0) <= fifo_full_140097944128592(0);
        
        fifo_inputs_140097944128648(0) <= outputs_140097944128592(0);
        outputs_full_140097944128592(0) <= fifo_full_140097944128648(0);
        
        fifo_inputs_140097944128704(0) <= outputs_140097944128648(0);
        outputs_full_140097944128648(0) <= fifo_full_140097944128704(0);
        
        fifo_inputs_140097944128760(0) <= outputs_140097944128704(0);
        outputs_full_140097944128704(0) <= fifo_full_140097944128760(0);
        
        fifo_inputs_140097944128816(0) <= outputs_140097944128760(0);
        outputs_full_140097944128760(0) <= fifo_full_140097944128816(0);
        
        fifo_inputs_140097944128872(0) <= outputs_140097944128816(0);
        outputs_full_140097944128816(0) <= fifo_full_140097944128872(0);
        
        fifo_inputs_140097944128928(0) <= outputs_140097944128872(0);
        outputs_full_140097944128872(0) <= fifo_full_140097944128928(0);
        
        fifo_inputs_140097944128984(0) <= outputs_140097944128928(0);
        outputs_full_140097944128928(0) <= fifo_full_140097944128984(0);
        
        fifo_inputs_140097944129040(0) <= outputs_140097944128984(0);
        outputs_full_140097944128984(0) <= fifo_full_140097944129040(0);
        
        fifo_inputs_140097944129096(0) <= outputs_140097944129040(0);
        outputs_full_140097944129040(0) <= fifo_full_140097944129096(0);
        
        fifo_inputs_140097944129152(0) <= outputs_140097944129096(0);
        outputs_full_140097944129096(0) <= fifo_full_140097944129152(0);
        
        fifo_inputs_140097944129208(0) <= outputs_140097944129152(0);
        outputs_full_140097944129152(0) <= fifo_full_140097944129208(0);
        
        fifo_inputs_140097944129264(0) <= outputs_140097944129208(0);
        outputs_full_140097944129208(0) <= fifo_full_140097944129264(0);
        
        fifo_inputs_140097944129320(0) <= outputs_140097944129264(0);
        outputs_full_140097944129264(0) <= fifo_full_140097944129320(0);
        
        fifo_inputs_140097944129376(0) <= outputs_140097944129320(0);
        outputs_full_140097944129320(0) <= fifo_full_140097944129376(0);
        
        fifo_inputs_140097944129432(0) <= outputs_140097944129376(0);
        outputs_full_140097944129376(0) <= fifo_full_140097944129432(0);
        
        fifo_inputs_140097944129488(0) <= outputs_140097944129432(0);
        outputs_full_140097944129432(0) <= fifo_full_140097944129488(0);
        
        fifo_inputs_140097944141896(0) <= outputs_140097944129488(0);
        outputs_full_140097944129488(0) <= fifo_full_140097944141896(0);
        
        fifo_inputs_140097944141952(0) <= outputs_140097944141896(0);
        outputs_full_140097944141896(0) <= fifo_full_140097944141952(0);
        
        fifo_inputs_140097944142008(0) <= outputs_140097944141952(0);
        outputs_full_140097944141952(0) <= fifo_full_140097944142008(0);
        
        fifo_inputs_140097944142064(0) <= outputs_140097944142008(0);
        outputs_full_140097944142008(0) <= fifo_full_140097944142064(0);
        
        fifo_inputs_140097944142120(0) <= outputs_140097944142064(0);
        outputs_full_140097944142064(0) <= fifo_full_140097944142120(0);
        
        fifo_inputs_140097944142176(0) <= outputs_140097944142120(0);
        outputs_full_140097944142120(0) <= fifo_full_140097944142176(0);
        
        fifo_inputs_140097944142232(0) <= outputs_140097944142176(0);
        outputs_full_140097944142176(0) <= fifo_full_140097944142232(0);
        
        fifo_inputs_140097944142288(0) <= outputs_140097944142232(0);
        outputs_full_140097944142232(0) <= fifo_full_140097944142288(0);
        
        fifo_inputs_140097944142344(0) <= outputs_140097944142288(0);
        outputs_full_140097944142288(0) <= fifo_full_140097944142344(0);
        
        fifo_inputs_140097944142400(0) <= outputs_140097944142344(0);
        outputs_full_140097944142344(0) <= fifo_full_140097944142400(0);
        
        fifo_inputs_140097944142456(0) <= outputs_140097944142400(0);
        outputs_full_140097944142400(0) <= fifo_full_140097944142456(0);
        
        fifo_inputs_140097944142512(0) <= outputs_140097944142456(0);
        outputs_full_140097944142456(0) <= fifo_full_140097944142512(0);
        
        fifo_inputs_140097944142568(0) <= outputs_140097944142512(0);
        outputs_full_140097944142512(0) <= fifo_full_140097944142568(0);
        
        fifo_inputs_140097944142624(0) <= outputs_140097944142568(0);
        outputs_full_140097944142568(0) <= fifo_full_140097944142624(0);
        
        fifo_inputs_140097944142680(0) <= outputs_140097944142624(0);
        outputs_full_140097944142624(0) <= fifo_full_140097944142680(0);
        
        fifo_inputs_140097944142736(0) <= outputs_140097944142680(0);
        outputs_full_140097944142680(0) <= fifo_full_140097944142736(0);
        
        fifo_inputs_140097944142792(0) <= outputs_140097944142736(0);
        outputs_full_140097944142736(0) <= fifo_full_140097944142792(0);
        
        fifo_inputs_140097944142848(0) <= outputs_140097944142792(0);
        outputs_full_140097944142792(0) <= fifo_full_140097944142848(0);
        
        fifo_inputs_140097944142904(0) <= outputs_140097944142848(0);
        outputs_full_140097944142848(0) <= fifo_full_140097944142904(0);
        
        fifo_inputs_140097944142960(0) <= outputs_140097944142904(0);
        outputs_full_140097944142904(0) <= fifo_full_140097944142960(0);
        
        fifo_inputs_140097944143016(0) <= outputs_140097944142960(0);
        outputs_full_140097944142960(0) <= fifo_full_140097944143016(0);
        
        fifo_inputs_140097944143072(0) <= outputs_140097944143016(0);
        outputs_full_140097944143016(0) <= fifo_full_140097944143072(0);
        
        fifo_inputs_140097944143128(0) <= outputs_140097944143072(0);
        outputs_full_140097944143072(0) <= fifo_full_140097944143128(0);
        
        fifo_inputs_140097944143184(0) <= outputs_140097944143128(0);
        outputs_full_140097944143128(0) <= fifo_full_140097944143184(0);
        
        fifo_inputs_140097944143240(0) <= outputs_140097944143184(0);
        outputs_full_140097944143184(0) <= fifo_full_140097944143240(0);
        
        fifo_inputs_140097944143296(0) <= outputs_140097944143240(0);
        outputs_full_140097944143240(0) <= fifo_full_140097944143296(0);
        
        fifo_inputs_140097944143352(0) <= outputs_140097944143296(0);
        outputs_full_140097944143296(0) <= fifo_full_140097944143352(0);
        
        fifo_inputs_140097944143408(0) <= outputs_140097944143352(0);
        outputs_full_140097944143352(0) <= fifo_full_140097944143408(0);
        
        fifo_inputs_140097944143464(0) <= outputs_140097944143408(0);
        outputs_full_140097944143408(0) <= fifo_full_140097944143464(0);
        
        fifo_inputs_140097944143520(0) <= outputs_140097944143464(0);
        outputs_full_140097944143464(0) <= fifo_full_140097944143520(0);
        
        fifo_inputs_140097944143576(0) <= outputs_140097944143520(0);
        outputs_full_140097944143520(0) <= fifo_full_140097944143576(0);
        
        fifo_inputs_140097944143632(0) <= outputs_140097944143576(0);
        outputs_full_140097944143576(0) <= fifo_full_140097944143632(0);
        
        fifo_inputs_140097944143688(0) <= outputs_140097944143632(0);
        outputs_full_140097944143632(0) <= fifo_full_140097944143688(0);
        
        fifo_inputs_140097944143744(0) <= outputs_140097944143688(0);
        outputs_full_140097944143688(0) <= fifo_full_140097944143744(0);
        
        fifo_inputs_140097944143800(0) <= outputs_140097944143744(0);
        outputs_full_140097944143744(0) <= fifo_full_140097944143800(0);
        
        fifo_inputs_140097944143856(0) <= outputs_140097944143800(0);
        outputs_full_140097944143800(0) <= fifo_full_140097944143856(0);
        
        fifo_inputs_140097944143912(0) <= outputs_140097944143856(0);
        outputs_full_140097944143856(0) <= fifo_full_140097944143912(0);
        
        fifo_inputs_140097944143968(0) <= outputs_140097944143912(0);
        outputs_full_140097944143912(0) <= fifo_full_140097944143968(0);
        
        fifo_inputs_140097944144024(0) <= outputs_140097944143968(0);
        outputs_full_140097944143968(0) <= fifo_full_140097944144024(0);
        
        fifo_inputs_140097944144080(0) <= outputs_140097944144024(0);
        outputs_full_140097944144024(0) <= fifo_full_140097944144080(0);
        
        fifo_inputs_140097944144136(0) <= outputs_140097944144080(0);
        outputs_full_140097944144080(0) <= fifo_full_140097944144136(0);
        
        fifo_inputs_140097944144192(0) <= outputs_140097944144136(0);
        outputs_full_140097944144136(0) <= fifo_full_140097944144192(0);
        
        fifo_inputs_140097944144248(0) <= outputs_140097944144192(0);
        outputs_full_140097944144192(0) <= fifo_full_140097944144248(0);
        
        fifo_inputs_140097944144304(0) <= outputs_140097944144248(0);
        outputs_full_140097944144248(0) <= fifo_full_140097944144304(0);
        
        fifo_inputs_140097944144360(0) <= outputs_140097944144304(0);
        outputs_full_140097944144304(0) <= fifo_full_140097944144360(0);
        
        fifo_inputs_140097944144416(0) <= outputs_140097944144360(0);
        outputs_full_140097944144360(0) <= fifo_full_140097944144416(0);
        
        fifo_inputs_140097944144472(0) <= outputs_140097944144416(0);
        outputs_full_140097944144416(0) <= fifo_full_140097944144472(0);
        
        fifo_inputs_140097944144528(0) <= outputs_140097944144472(0);
        outputs_full_140097944144472(0) <= fifo_full_140097944144528(0);
        
        fifo_inputs_140097944144584(0) <= outputs_140097944144528(0);
        outputs_full_140097944144528(0) <= fifo_full_140097944144584(0);
        
        fifo_inputs_140097944144640(0) <= outputs_140097944144584(0);
        outputs_full_140097944144584(0) <= fifo_full_140097944144640(0);
        
        fifo_inputs_140097944144696(0) <= outputs_140097944144640(0);
        outputs_full_140097944144640(0) <= fifo_full_140097944144696(0);
        
        fifo_inputs_140097944144752(0) <= outputs_140097944144696(0);
        outputs_full_140097944144696(0) <= fifo_full_140097944144752(0);
        
        fifo_inputs_140097944144808(0) <= outputs_140097944144752(0);
        outputs_full_140097944144752(0) <= fifo_full_140097944144808(0);
        
        fifo_inputs_140097944144864(0) <= outputs_140097944144808(0);
        outputs_full_140097944144808(0) <= fifo_full_140097944144864(0);
        
        fifo_inputs_140097944144920(0) <= outputs_140097944144864(0);
        outputs_full_140097944144864(0) <= fifo_full_140097944144920(0);
        
        fifo_inputs_140097944144976(0) <= outputs_140097944144920(0);
        outputs_full_140097944144920(0) <= fifo_full_140097944144976(0);
        
        fifo_inputs_140097944145032(0) <= outputs_140097944144976(0);
        outputs_full_140097944144976(0) <= fifo_full_140097944145032(0);
        
        fifo_inputs_140097944145088(0) <= outputs_140097944145032(0);
        outputs_full_140097944145032(0) <= fifo_full_140097944145088(0);
        
        fifo_inputs_140097944145144(0) <= outputs_140097944145088(0);
        outputs_full_140097944145088(0) <= fifo_full_140097944145144(0);
        
        fifo_inputs_140097944145200(0) <= outputs_140097944145144(0);
        outputs_full_140097944145144(0) <= fifo_full_140097944145200(0);
        
        fifo_inputs_140097944145256(0) <= outputs_140097944145200(0);
        outputs_full_140097944145200(0) <= fifo_full_140097944145256(0);
        
        fifo_inputs_140097944145312(0) <= outputs_140097944145256(0);
        outputs_full_140097944145256(0) <= fifo_full_140097944145312(0);
        
        fifo_inputs_140097944145368(0) <= outputs_140097944145312(0);
        outputs_full_140097944145312(0) <= fifo_full_140097944145368(0);
        
        fifo_inputs_140097944145424(0) <= outputs_140097944145368(0);
        outputs_full_140097944145368(0) <= fifo_full_140097944145424(0);
        
        fifo_inputs_140097944145480(0) <= outputs_140097944145424(0);
        outputs_full_140097944145424(0) <= fifo_full_140097944145480(0);
        
        fifo_inputs_140097944145536(0) <= outputs_140097944145480(0);
        outputs_full_140097944145480(0) <= fifo_full_140097944145536(0);
        
        fifo_inputs_140097944145592(0) <= outputs_140097944145536(0);
        outputs_full_140097944145536(0) <= fifo_full_140097944145592(0);
        
        fifo_inputs_140097944145648(0) <= outputs_140097944145592(0);
        outputs_full_140097944145592(0) <= fifo_full_140097944145648(0);
        
        fifo_inputs_140097944145704(0) <= outputs_140097944145648(0);
        outputs_full_140097944145648(0) <= fifo_full_140097944145704(0);
        
        fifo_inputs_140097944145760(0) <= outputs_140097944145704(0);
        outputs_full_140097944145704(0) <= fifo_full_140097944145760(0);
        
        fifo_inputs_140097944145816(0) <= outputs_140097944145760(0);
        outputs_full_140097944145760(0) <= fifo_full_140097944145816(0);
        
        fifo_inputs_140097944145872(0) <= outputs_140097944145816(0);
        outputs_full_140097944145816(0) <= fifo_full_140097944145872(0);
        
        fifo_inputs_140097944154184(0) <= outputs_140097944145872(0);
        outputs_full_140097944145872(0) <= fifo_full_140097944154184(0);
        
        fifo_inputs_140097944154240(0) <= outputs_140097944154184(0);
        outputs_full_140097944154184(0) <= fifo_full_140097944154240(0);
        
        fifo_inputs_140097944154296(0) <= outputs_140097944154240(0);
        outputs_full_140097944154240(0) <= fifo_full_140097944154296(0);
        
        fifo_inputs_140097944154352(0) <= outputs_140097944154296(0);
        outputs_full_140097944154296(0) <= fifo_full_140097944154352(0);
        
        fifo_inputs_140097944154408(0) <= outputs_140097944154352(0);
        outputs_full_140097944154352(0) <= fifo_full_140097944154408(0);
        
        fifo_inputs_140097944154464(0) <= outputs_140097944154408(0);
        outputs_full_140097944154408(0) <= fifo_full_140097944154464(0);
        
        fifo_inputs_140097944154520(0) <= outputs_140097944154464(0);
        outputs_full_140097944154464(0) <= fifo_full_140097944154520(0);
        
        fifo_inputs_140097944154576(0) <= outputs_140097944154520(0);
        outputs_full_140097944154520(0) <= fifo_full_140097944154576(0);
        
        fifo_inputs_140097944154632(0) <= outputs_140097944154576(0);
        outputs_full_140097944154576(0) <= fifo_full_140097944154632(0);
        
        fifo_inputs_140097944154688(0) <= outputs_140097944154632(0);
        outputs_full_140097944154632(0) <= fifo_full_140097944154688(0);
        
        fifo_inputs_140097944154744(0) <= outputs_140097944154688(0);
        outputs_full_140097944154688(0) <= fifo_full_140097944154744(0);
        
        fifo_inputs_140097944154800(0) <= outputs_140097944154744(0);
        outputs_full_140097944154744(0) <= fifo_full_140097944154800(0);
        
        fifo_inputs_140097944154856(0) <= outputs_140097944154800(0);
        outputs_full_140097944154800(0) <= fifo_full_140097944154856(0);
        
        fifo_inputs_140097944154912(0) <= outputs_140097944154856(0);
        outputs_full_140097944154856(0) <= fifo_full_140097944154912(0);
        
        fifo_inputs_140097944154968(0) <= outputs_140097944154912(0);
        outputs_full_140097944154912(0) <= fifo_full_140097944154968(0);
        
        fifo_inputs_140097944155024(0) <= outputs_140097944154968(0);
        outputs_full_140097944154968(0) <= fifo_full_140097944155024(0);
        
        fifo_inputs_140097944155080(0) <= outputs_140097944155024(0);
        outputs_full_140097944155024(0) <= fifo_full_140097944155080(0);
        
        fifo_inputs_140097944155136(0) <= outputs_140097944155080(0);
        outputs_full_140097944155080(0) <= fifo_full_140097944155136(0);
        
        fifo_inputs_140097944155192(0) <= outputs_140097944155136(0);
        outputs_full_140097944155136(0) <= fifo_full_140097944155192(0);
        
        fifo_inputs_140097944155248(0) <= outputs_140097944155192(0);
        outputs_full_140097944155192(0) <= fifo_full_140097944155248(0);
        
        fifo_inputs_140097944155304(0) <= outputs_140097944155248(0);
        outputs_full_140097944155248(0) <= fifo_full_140097944155304(0);
        
        fifo_inputs_140097944155360(0) <= outputs_140097944155304(0);
        outputs_full_140097944155304(0) <= fifo_full_140097944155360(0);
        
        fifo_inputs_140097944155416(0) <= outputs_140097944155360(0);
        outputs_full_140097944155360(0) <= fifo_full_140097944155416(0);
        
        fifo_inputs_140097944155472(0) <= outputs_140097944155416(0);
        outputs_full_140097944155416(0) <= fifo_full_140097944155472(0);
        
        fifo_inputs_140097944155528(0) <= outputs_140097944155472(0);
        outputs_full_140097944155472(0) <= fifo_full_140097944155528(0);
        
        fifo_inputs_140097944155584(0) <= outputs_140097944155528(0);
        outputs_full_140097944155528(0) <= fifo_full_140097944155584(0);
        
        fifo_inputs_140097944155640(0) <= outputs_140097944155584(0);
        outputs_full_140097944155584(0) <= fifo_full_140097944155640(0);
        
        fifo_inputs_140097944155696(0) <= outputs_140097944155640(0);
        outputs_full_140097944155640(0) <= fifo_full_140097944155696(0);
        
        fifo_inputs_140097944155752(0) <= outputs_140097944155696(0);
        outputs_full_140097944155696(0) <= fifo_full_140097944155752(0);
        
        fifo_inputs_140097944155808(0) <= outputs_140097944155752(0);
        outputs_full_140097944155752(0) <= fifo_full_140097944155808(0);
        
        fifo_inputs_140097944155864(0) <= outputs_140097944155808(0);
        outputs_full_140097944155808(0) <= fifo_full_140097944155864(0);
        
        fifo_inputs_140097944155920(0) <= outputs_140097944155864(0);
        outputs_full_140097944155864(0) <= fifo_full_140097944155920(0);
        
        fifo_inputs_140097944155976(0) <= outputs_140097944155920(0);
        outputs_full_140097944155920(0) <= fifo_full_140097944155976(0);
        
        fifo_inputs_140097944156032(0) <= outputs_140097944155976(0);
        outputs_full_140097944155976(0) <= fifo_full_140097944156032(0);
        
        fifo_inputs_140097944156088(0) <= outputs_140097944156032(0);
        outputs_full_140097944156032(0) <= fifo_full_140097944156088(0);
        
        fifo_inputs_140097944156144(0) <= outputs_140097944156088(0);
        outputs_full_140097944156088(0) <= fifo_full_140097944156144(0);
        
        fifo_inputs_140097944156200(0) <= outputs_140097944156144(0);
        outputs_full_140097944156144(0) <= fifo_full_140097944156200(0);
        
        fifo_inputs_140097944156256(0) <= outputs_140097944156200(0);
        outputs_full_140097944156200(0) <= fifo_full_140097944156256(0);
        
        fifo_inputs_140097944156312(0) <= outputs_140097944156256(0);
        outputs_full_140097944156256(0) <= fifo_full_140097944156312(0);
        
        fifo_inputs_140097944156368(0) <= outputs_140097944156312(0);
        outputs_full_140097944156312(0) <= fifo_full_140097944156368(0);
        
        fifo_inputs_140097944156424(0) <= outputs_140097944156368(0);
        outputs_full_140097944156368(0) <= fifo_full_140097944156424(0);
        
        fifo_inputs_140097944156480(0) <= outputs_140097944156424(0);
        outputs_full_140097944156424(0) <= fifo_full_140097944156480(0);
        
        fifo_inputs_140097944156536(0) <= outputs_140097944156480(0);
        outputs_full_140097944156480(0) <= fifo_full_140097944156536(0);
        
        fifo_inputs_140097944156592(0) <= outputs_140097944156536(0);
        outputs_full_140097944156536(0) <= fifo_full_140097944156592(0);
        
        fifo_inputs_140097944156648(0) <= outputs_140097944156592(0);
        outputs_full_140097944156592(0) <= fifo_full_140097944156648(0);
        
        fifo_inputs_140097944156704(0) <= outputs_140097944156648(0);
        outputs_full_140097944156648(0) <= fifo_full_140097944156704(0);
        
        fifo_inputs_140097944156760(0) <= outputs_140097944156704(0);
        outputs_full_140097944156704(0) <= fifo_full_140097944156760(0);
        
        fifo_inputs_140097944156816(0) <= outputs_140097944156760(0);
        outputs_full_140097944156760(0) <= fifo_full_140097944156816(0);
        
        fifo_inputs_140097944156872(0) <= outputs_140097944156816(0);
        outputs_full_140097944156816(0) <= fifo_full_140097944156872(0);
        
        fifo_inputs_140097944156928(0) <= outputs_140097944156872(0);
        outputs_full_140097944156872(0) <= fifo_full_140097944156928(0);
        
        fifo_inputs_140097944156984(0) <= outputs_140097944156928(0);
        outputs_full_140097944156928(0) <= fifo_full_140097944156984(0);
        
        fifo_inputs_140097944157040(0) <= outputs_140097944156984(0);
        outputs_full_140097944156984(0) <= fifo_full_140097944157040(0);
        
        fifo_inputs_140097944157096(0) <= outputs_140097944157040(0);
        outputs_full_140097944157040(0) <= fifo_full_140097944157096(0);
        
        fifo_inputs_140097944157152(0) <= outputs_140097944157096(0);
        outputs_full_140097944157096(0) <= fifo_full_140097944157152(0);
        
        fifo_inputs_140097944157208(0) <= outputs_140097944157152(0);
        outputs_full_140097944157152(0) <= fifo_full_140097944157208(0);
        
        fifo_inputs_140097944157264(0) <= outputs_140097944157208(0);
        outputs_full_140097944157208(0) <= fifo_full_140097944157264(0);
        
        fifo_inputs_140097944157320(0) <= outputs_140097944157264(0);
        outputs_full_140097944157264(0) <= fifo_full_140097944157320(0);
        
        fifo_inputs_140097944157376(0) <= outputs_140097944157320(0);
        outputs_full_140097944157320(0) <= fifo_full_140097944157376(0);
        
        fifo_inputs_140097944157432(0) <= outputs_140097944157376(0);
        outputs_full_140097944157376(0) <= fifo_full_140097944157432(0);
        
        fifo_inputs_140097944157488(0) <= outputs_140097944157432(0);
        outputs_full_140097944157432(0) <= fifo_full_140097944157488(0);
        
        fifo_inputs_140097944157544(0) <= outputs_140097944157488(0);
        outputs_full_140097944157488(0) <= fifo_full_140097944157544(0);
        
        fifo_inputs_140097944157600(0) <= outputs_140097944157544(0);
        outputs_full_140097944157544(0) <= fifo_full_140097944157600(0);
        
        fifo_inputs_140097944157656(0) <= outputs_140097944157600(0);
        outputs_full_140097944157600(0) <= fifo_full_140097944157656(0);
        
        fifo_inputs_140097944157712(0) <= outputs_140097944157656(0);
        outputs_full_140097944157656(0) <= fifo_full_140097944157712(0);
        
        fifo_inputs_140097944157768(0) <= outputs_140097944157712(0);
        outputs_full_140097944157712(0) <= fifo_full_140097944157768(0);
        
        fifo_inputs_140097944157824(0) <= outputs_140097944157768(0);
        outputs_full_140097944157768(0) <= fifo_full_140097944157824(0);
        
        fifo_inputs_140097944157880(0) <= outputs_140097944157824(0);
        outputs_full_140097944157824(0) <= fifo_full_140097944157880(0);
        
        fifo_inputs_140097944157936(0) <= outputs_140097944157880(0);
        outputs_full_140097944157880(0) <= fifo_full_140097944157936(0);
        
        fifo_inputs_140097944157992(0) <= outputs_140097944157936(0);
        outputs_full_140097944157936(0) <= fifo_full_140097944157992(0);
        
        fifo_inputs_140097944158048(0) <= outputs_140097944157992(0);
        outputs_full_140097944157992(0) <= fifo_full_140097944158048(0);
        
        fifo_inputs_140097944158104(0) <= outputs_140097944158048(0);
        outputs_full_140097944158048(0) <= fifo_full_140097944158104(0);
        
        fifo_inputs_140097944158160(0) <= outputs_140097944158104(0);
        outputs_full_140097944158104(0) <= fifo_full_140097944158160(0);
        
        fifo_inputs_140097944166472(0) <= outputs_140097944158160(0);
        outputs_full_140097944158160(0) <= fifo_full_140097944166472(0);
        
        fifo_inputs_140097944166528(0) <= outputs_140097944166472(0);
        outputs_full_140097944166472(0) <= fifo_full_140097944166528(0);
        
        fifo_inputs_140097944166584(0) <= outputs_140097944166528(0);
        outputs_full_140097944166528(0) <= fifo_full_140097944166584(0);
        
        fifo_inputs_140097944166640(0) <= outputs_140097944166584(0);
        outputs_full_140097944166584(0) <= fifo_full_140097944166640(0);
        
        fifo_inputs_140097944166696(0) <= outputs_140097944166640(0);
        outputs_full_140097944166640(0) <= fifo_full_140097944166696(0);
        
        fifo_inputs_140097944166752(0) <= outputs_140097944166696(0);
        outputs_full_140097944166696(0) <= fifo_full_140097944166752(0);
        
        fifo_inputs_140097944166808(0) <= outputs_140097944166752(0);
        outputs_full_140097944166752(0) <= fifo_full_140097944166808(0);
        
        fifo_inputs_140097944166864(0) <= outputs_140097944166808(0);
        outputs_full_140097944166808(0) <= fifo_full_140097944166864(0);
        
        fifo_inputs_140097944166920(0) <= outputs_140097944166864(0);
        outputs_full_140097944166864(0) <= fifo_full_140097944166920(0);
        
        fifo_inputs_140097944166976(0) <= outputs_140097944166920(0);
        outputs_full_140097944166920(0) <= fifo_full_140097944166976(0);
        
        fifo_inputs_140097944167032(0) <= outputs_140097944166976(0);
        outputs_full_140097944166976(0) <= fifo_full_140097944167032(0);
        
        fifo_inputs_140097944167088(0) <= outputs_140097944167032(0);
        outputs_full_140097944167032(0) <= fifo_full_140097944167088(0);
        
        fifo_inputs_140097944167144(0) <= outputs_140097944167088(0);
        outputs_full_140097944167088(0) <= fifo_full_140097944167144(0);
        
        fifo_inputs_140097944167200(0) <= outputs_140097944167144(0);
        outputs_full_140097944167144(0) <= fifo_full_140097944167200(0);
        
        fifo_inputs_140097944167256(0) <= outputs_140097944167200(0);
        outputs_full_140097944167200(0) <= fifo_full_140097944167256(0);
        
        fifo_inputs_140097944167312(0) <= outputs_140097944167256(0);
        outputs_full_140097944167256(0) <= fifo_full_140097944167312(0);
        
        fifo_inputs_140097944167368(0) <= outputs_140097944167312(0);
        outputs_full_140097944167312(0) <= fifo_full_140097944167368(0);
        
        fifo_inputs_140097944167424(0) <= outputs_140097944167368(0);
        outputs_full_140097944167368(0) <= fifo_full_140097944167424(0);
        
        fifo_inputs_140097944167480(0) <= outputs_140097944167424(0);
        outputs_full_140097944167424(0) <= fifo_full_140097944167480(0);
        
        fifo_inputs_140097944167536(0) <= outputs_140097944167480(0);
        outputs_full_140097944167480(0) <= fifo_full_140097944167536(0);
        
        fifo_inputs_140097944167592(0) <= outputs_140097944167536(0);
        outputs_full_140097944167536(0) <= fifo_full_140097944167592(0);
        
        fifo_inputs_140097944167648(0) <= outputs_140097944167592(0);
        outputs_full_140097944167592(0) <= fifo_full_140097944167648(0);
        
        fifo_inputs_140097944167704(0) <= outputs_140097944167648(0);
        outputs_full_140097944167648(0) <= fifo_full_140097944167704(0);
        
        fifo_inputs_140097944167760(0) <= outputs_140097944167704(0);
        outputs_full_140097944167704(0) <= fifo_full_140097944167760(0);
        
        fifo_inputs_140097944167816(0) <= outputs_140097944167760(0);
        outputs_full_140097944167760(0) <= fifo_full_140097944167816(0);
        
        fifo_inputs_140097944167872(0) <= outputs_140097944167816(0);
        outputs_full_140097944167816(0) <= fifo_full_140097944167872(0);
        
        fifo_inputs_140097944167928(0) <= outputs_140097944167872(0);
        outputs_full_140097944167872(0) <= fifo_full_140097944167928(0);
        
        fifo_inputs_140097944167984(0) <= outputs_140097944167928(0);
        outputs_full_140097944167928(0) <= fifo_full_140097944167984(0);
        
        fifo_inputs_140097944168040(0) <= outputs_140097944167984(0);
        outputs_full_140097944167984(0) <= fifo_full_140097944168040(0);
        
        fifo_inputs_140097944168096(0) <= outputs_140097944168040(0);
        outputs_full_140097944168040(0) <= fifo_full_140097944168096(0);
        
        fifo_inputs_140097944168152(0) <= outputs_140097944168096(0);
        outputs_full_140097944168096(0) <= fifo_full_140097944168152(0);
        
        fifo_inputs_140097944168208(0) <= outputs_140097944168152(0);
        outputs_full_140097944168152(0) <= fifo_full_140097944168208(0);
        
        fifo_inputs_140097944168264(0) <= outputs_140097944168208(0);
        outputs_full_140097944168208(0) <= fifo_full_140097944168264(0);
        
        fifo_inputs_140097944168320(0) <= outputs_140097944168264(0);
        outputs_full_140097944168264(0) <= fifo_full_140097944168320(0);
        
        fifo_inputs_140097944168376(0) <= outputs_140097944168320(0);
        outputs_full_140097944168320(0) <= fifo_full_140097944168376(0);
        
        fifo_inputs_140097944168432(0) <= outputs_140097944168376(0);
        outputs_full_140097944168376(0) <= fifo_full_140097944168432(0);
        
        fifo_inputs_140097944168488(0) <= outputs_140097944168432(0);
        outputs_full_140097944168432(0) <= fifo_full_140097944168488(0);
        
        fifo_inputs_140097944168544(0) <= outputs_140097944168488(0);
        outputs_full_140097944168488(0) <= fifo_full_140097944168544(0);
        
        fifo_inputs_140097944168600(0) <= outputs_140097944168544(0);
        outputs_full_140097944168544(0) <= fifo_full_140097944168600(0);
        
        fifo_inputs_140097944168656(0) <= outputs_140097944168600(0);
        outputs_full_140097944168600(0) <= fifo_full_140097944168656(0);
        
        fifo_inputs_140097944168712(0) <= outputs_140097944168656(0);
        outputs_full_140097944168656(0) <= fifo_full_140097944168712(0);
        
        fifo_inputs_140097944168768(0) <= outputs_140097944168712(0);
        outputs_full_140097944168712(0) <= fifo_full_140097944168768(0);
        
        fifo_inputs_140097944168824(0) <= outputs_140097944168768(0);
        outputs_full_140097944168768(0) <= fifo_full_140097944168824(0);
        
        fifo_inputs_140097944168880(0) <= outputs_140097944168824(0);
        outputs_full_140097944168824(0) <= fifo_full_140097944168880(0);
        
        fifo_inputs_140097944168936(0) <= outputs_140097944168880(0);
        outputs_full_140097944168880(0) <= fifo_full_140097944168936(0);
        
        fifo_inputs_140097944168992(0) <= outputs_140097944168936(0);
        outputs_full_140097944168936(0) <= fifo_full_140097944168992(0);
        
        fifo_inputs_140097944169048(0) <= outputs_140097944168992(0);
        outputs_full_140097944168992(0) <= fifo_full_140097944169048(0);
        
        fifo_inputs_140097944169104(0) <= outputs_140097944169048(0);
        outputs_full_140097944169048(0) <= fifo_full_140097944169104(0);
        
        fifo_inputs_140097944169160(0) <= outputs_140097944169104(0);
        outputs_full_140097944169104(0) <= fifo_full_140097944169160(0);
        
        fifo_inputs_140097944169216(0) <= outputs_140097944169160(0);
        outputs_full_140097944169160(0) <= fifo_full_140097944169216(0);
        
        fifo_inputs_140097944169272(0) <= outputs_140097944169216(0);
        outputs_full_140097944169216(0) <= fifo_full_140097944169272(0);
        
        fifo_inputs_140097944169328(0) <= outputs_140097944169272(0);
        outputs_full_140097944169272(0) <= fifo_full_140097944169328(0);
        
        fifo_inputs_140097944169384(0) <= outputs_140097944169328(0);
        outputs_full_140097944169328(0) <= fifo_full_140097944169384(0);
        
        fifo_inputs_140097944169440(0) <= outputs_140097944169384(0);
        outputs_full_140097944169384(0) <= fifo_full_140097944169440(0);
        
        fifo_inputs_140097944169496(0) <= outputs_140097944169440(0);
        outputs_full_140097944169440(0) <= fifo_full_140097944169496(0);
        
        fifo_inputs_140097944169552(0) <= outputs_140097944169496(0);
        outputs_full_140097944169496(0) <= fifo_full_140097944169552(0);
        
        fifo_inputs_140097944169608(0) <= outputs_140097944169552(0);
        outputs_full_140097944169552(0) <= fifo_full_140097944169608(0);
        
        fifo_inputs_140097944169664(0) <= outputs_140097944169608(0);
        outputs_full_140097944169608(0) <= fifo_full_140097944169664(0);
        
        fifo_inputs_140097944169720(0) <= outputs_140097944169664(0);
        outputs_full_140097944169664(0) <= fifo_full_140097944169720(0);
        
        fifo_inputs_140097944169776(0) <= outputs_140097944169720(0);
        outputs_full_140097944169720(0) <= fifo_full_140097944169776(0);
        
        fifo_inputs_140097944169832(0) <= outputs_140097944169776(0);
        outputs_full_140097944169776(0) <= fifo_full_140097944169832(0);
        
        fifo_inputs_140097944169888(0) <= outputs_140097944169832(0);
        outputs_full_140097944169832(0) <= fifo_full_140097944169888(0);
        
        fifo_inputs_140097944169944(0) <= outputs_140097944169888(0);
        outputs_full_140097944169888(0) <= fifo_full_140097944169944(0);
        
        fifo_inputs_140097944170000(0) <= outputs_140097944169944(0);
        outputs_full_140097944169944(0) <= fifo_full_140097944170000(0);
        
        fifo_inputs_140097944170056(0) <= outputs_140097944170000(0);
        outputs_full_140097944170000(0) <= fifo_full_140097944170056(0);
        
        fifo_inputs_140097944170112(0) <= outputs_140097944170056(0);
        outputs_full_140097944170056(0) <= fifo_full_140097944170112(0);
        
        fifo_inputs_140097944170168(0) <= outputs_140097944170112(0);
        outputs_full_140097944170112(0) <= fifo_full_140097944170168(0);
        
        fifo_inputs_140097944170224(0) <= outputs_140097944170168(0);
        outputs_full_140097944170168(0) <= fifo_full_140097944170224(0);
        
        fifo_inputs_140097944170280(0) <= outputs_140097944170224(0);
        outputs_full_140097944170224(0) <= fifo_full_140097944170280(0);
        
        fifo_inputs_140097944170336(0) <= outputs_140097944170280(0);
        outputs_full_140097944170280(0) <= fifo_full_140097944170336(0);
        
        fifo_inputs_140097944170392(0) <= outputs_140097944170336(0);
        outputs_full_140097944170336(0) <= fifo_full_140097944170392(0);
        
        fifo_inputs_140097944170448(0) <= outputs_140097944170392(0);
        outputs_full_140097944170392(0) <= fifo_full_140097944170448(0);
        
        fifo_inputs_140097941516360(0) <= outputs_140097944170448(0);
        outputs_full_140097944170448(0) <= fifo_full_140097941516360(0);
        
        fifo_inputs_140097941516416(0) <= outputs_140097941516360(0);
        outputs_full_140097941516360(0) <= fifo_full_140097941516416(0);
        
        fifo_inputs_140097941516472(0) <= outputs_140097941516416(0);
        outputs_full_140097941516416(0) <= fifo_full_140097941516472(0);
        
        fifo_inputs_140097941516528(0) <= outputs_140097941516472(0);
        outputs_full_140097941516472(0) <= fifo_full_140097941516528(0);
        
        fifo_inputs_140097941516584(0) <= outputs_140097941516528(0);
        outputs_full_140097941516528(0) <= fifo_full_140097941516584(0);
        
        fifo_inputs_140097941516640(0) <= outputs_140097941516584(0);
        outputs_full_140097941516584(0) <= fifo_full_140097941516640(0);
        
        fifo_inputs_140097941516696(0) <= outputs_140097941516640(0);
        outputs_full_140097941516640(0) <= fifo_full_140097941516696(0);
        
        fifo_inputs_140097941516752(0) <= outputs_140097941516696(0);
        outputs_full_140097941516696(0) <= fifo_full_140097941516752(0);
        
        fifo_inputs_140097941516808(0) <= outputs_140097941516752(0);
        outputs_full_140097941516752(0) <= fifo_full_140097941516808(0);
        
        fifo_inputs_140097941516864(0) <= outputs_140097941516808(0);
        outputs_full_140097941516808(0) <= fifo_full_140097941516864(0);
        
        fifo_inputs_140097941516920(0) <= outputs_140097941516864(0);
        outputs_full_140097941516864(0) <= fifo_full_140097941516920(0);
        
        fifo_inputs_140097941516976(0) <= outputs_140097941516920(0);
        outputs_full_140097941516920(0) <= fifo_full_140097941516976(0);
        
        fifo_inputs_140097941517032(0) <= outputs_140097941516976(0);
        outputs_full_140097941516976(0) <= fifo_full_140097941517032(0);
        
        fifo_inputs_140097941517088(0) <= outputs_140097941517032(0);
        outputs_full_140097941517032(0) <= fifo_full_140097941517088(0);
        
        fifo_inputs_140097941517144(0) <= outputs_140097941517088(0);
        outputs_full_140097941517088(0) <= fifo_full_140097941517144(0);
        
        fifo_inputs_140097941517200(0) <= outputs_140097941517144(0);
        outputs_full_140097941517144(0) <= fifo_full_140097941517200(0);
        
        fifo_inputs_140097941517256(0) <= outputs_140097941517200(0);
        outputs_full_140097941517200(0) <= fifo_full_140097941517256(0);
        
        fifo_inputs_140097941517312(0) <= outputs_140097941517256(0);
        outputs_full_140097941517256(0) <= fifo_full_140097941517312(0);
        
        fifo_inputs_140097941517368(0) <= outputs_140097941517312(0);
        outputs_full_140097941517312(0) <= fifo_full_140097941517368(0);
        
        fifo_inputs_140097941517424(0) <= outputs_140097941517368(0);
        outputs_full_140097941517368(0) <= fifo_full_140097941517424(0);
        
        fifo_inputs_140097941517480(0) <= outputs_140097941517424(0);
        outputs_full_140097941517424(0) <= fifo_full_140097941517480(0);
        
        fifo_inputs_140097941517536(0) <= outputs_140097941517480(0);
        outputs_full_140097941517480(0) <= fifo_full_140097941517536(0);
        
        fifo_inputs_140097941517592(0) <= outputs_140097941517536(0);
        outputs_full_140097941517536(0) <= fifo_full_140097941517592(0);
        
        fifo_inputs_140097941517648(0) <= outputs_140097941517592(0);
        outputs_full_140097941517592(0) <= fifo_full_140097941517648(0);
        
        fifo_inputs_140097941517704(0) <= outputs_140097941517648(0);
        outputs_full_140097941517648(0) <= fifo_full_140097941517704(0);
        
        fifo_inputs_140097941517760(0) <= outputs_140097941517704(0);
        outputs_full_140097941517704(0) <= fifo_full_140097941517760(0);
        
        fifo_inputs_140097941517816(0) <= outputs_140097941517760(0);
        outputs_full_140097941517760(0) <= fifo_full_140097941517816(0);
        
        fifo_inputs_140097941517872(0) <= outputs_140097941517816(0);
        outputs_full_140097941517816(0) <= fifo_full_140097941517872(0);
        
        fifo_inputs_140097941517928(0) <= outputs_140097941517872(0);
        outputs_full_140097941517872(0) <= fifo_full_140097941517928(0);
        
        fifo_inputs_140097941517984(0) <= outputs_140097941517928(0);
        outputs_full_140097941517928(0) <= fifo_full_140097941517984(0);
        
        fifo_inputs_140097941518040(0) <= outputs_140097941517984(0);
        outputs_full_140097941517984(0) <= fifo_full_140097941518040(0);
        
        fifo_inputs_140097941518096(0) <= outputs_140097941518040(0);
        outputs_full_140097941518040(0) <= fifo_full_140097941518096(0);
        
        fifo_inputs_140097941518152(0) <= outputs_140097941518096(0);
        outputs_full_140097941518096(0) <= fifo_full_140097941518152(0);
        
        fifo_inputs_140097941518208(0) <= outputs_140097941518152(0);
        outputs_full_140097941518152(0) <= fifo_full_140097941518208(0);
        
        fifo_inputs_140097941518264(0) <= outputs_140097941518208(0);
        outputs_full_140097941518208(0) <= fifo_full_140097941518264(0);
        
        fifo_inputs_140097941518320(0) <= outputs_140097941518264(0);
        outputs_full_140097941518264(0) <= fifo_full_140097941518320(0);
        
        fifo_inputs_140097941518376(0) <= outputs_140097941518320(0);
        outputs_full_140097941518320(0) <= fifo_full_140097941518376(0);
        
        fifo_inputs_140097941518432(0) <= outputs_140097941518376(0);
        outputs_full_140097941518376(0) <= fifo_full_140097941518432(0);
        
        fifo_inputs_140097941518488(0) <= outputs_140097941518432(0);
        outputs_full_140097941518432(0) <= fifo_full_140097941518488(0);
        
        fifo_inputs_140097941518544(0) <= outputs_140097941518488(0);
        outputs_full_140097941518488(0) <= fifo_full_140097941518544(0);
        
        fifo_inputs_140097941518600(0) <= outputs_140097941518544(0);
        outputs_full_140097941518544(0) <= fifo_full_140097941518600(0);
        
        fifo_inputs_140097941518656(0) <= outputs_140097941518600(0);
        outputs_full_140097941518600(0) <= fifo_full_140097941518656(0);
        
        fifo_inputs_140097941518712(0) <= outputs_140097941518656(0);
        outputs_full_140097941518656(0) <= fifo_full_140097941518712(0);
        
        fifo_inputs_140097941518768(0) <= outputs_140097941518712(0);
        outputs_full_140097941518712(0) <= fifo_full_140097941518768(0);
        
        fifo_inputs_140097941518824(0) <= outputs_140097941518768(0);
        outputs_full_140097941518768(0) <= fifo_full_140097941518824(0);
        
        fifo_inputs_140097941518880(0) <= outputs_140097941518824(0);
        outputs_full_140097941518824(0) <= fifo_full_140097941518880(0);
        
        fifo_inputs_140097941518936(0) <= outputs_140097941518880(0);
        outputs_full_140097941518880(0) <= fifo_full_140097941518936(0);
        
        fifo_inputs_140097941518992(0) <= outputs_140097941518936(0);
        outputs_full_140097941518936(0) <= fifo_full_140097941518992(0);
        
        fifo_inputs_140097941519048(0) <= outputs_140097941518992(0);
        outputs_full_140097941518992(0) <= fifo_full_140097941519048(0);
        
        fifo_inputs_140097941519104(0) <= outputs_140097941519048(0);
        outputs_full_140097941519048(0) <= fifo_full_140097941519104(0);
        
        fifo_inputs_140097941519160(0) <= outputs_140097941519104(0);
        outputs_full_140097941519104(0) <= fifo_full_140097941519160(0);
        
        fifo_inputs_140097941519216(0) <= outputs_140097941519160(0);
        outputs_full_140097941519160(0) <= fifo_full_140097941519216(0);
        
        fifo_inputs_140097941519272(0) <= outputs_140097941519216(0);
        outputs_full_140097941519216(0) <= fifo_full_140097941519272(0);
        
        fifo_inputs_140097941519328(0) <= outputs_140097941519272(0);
        outputs_full_140097941519272(0) <= fifo_full_140097941519328(0);
        
        fifo_inputs_140097941519384(0) <= outputs_140097941519328(0);
        outputs_full_140097941519328(0) <= fifo_full_140097941519384(0);
        
        fifo_inputs_140097941519440(0) <= outputs_140097941519384(0);
        outputs_full_140097941519384(0) <= fifo_full_140097941519440(0);
        
        fifo_inputs_140097941519496(0) <= outputs_140097941519440(0);
        outputs_full_140097941519440(0) <= fifo_full_140097941519496(0);
        
        fifo_inputs_140097941519552(0) <= outputs_140097941519496(0);
        outputs_full_140097941519496(0) <= fifo_full_140097941519552(0);
        
        fifo_inputs_140097941519608(0) <= outputs_140097941519552(0);
        outputs_full_140097941519552(0) <= fifo_full_140097941519608(0);
        
        fifo_inputs_140097941519664(0) <= outputs_140097941519608(0);
        outputs_full_140097941519608(0) <= fifo_full_140097941519664(0);
        
        fifo_inputs_140097941519720(0) <= outputs_140097941519664(0);
        outputs_full_140097941519664(0) <= fifo_full_140097941519720(0);
        
        fifo_inputs_140097941519776(0) <= outputs_140097941519720(0);
        outputs_full_140097941519720(0) <= fifo_full_140097941519776(0);
        
        fifo_inputs_140097941519832(0) <= outputs_140097941519776(0);
        outputs_full_140097941519776(0) <= fifo_full_140097941519832(0);
        
        fifo_inputs_140097941519888(0) <= outputs_140097941519832(0);
        outputs_full_140097941519832(0) <= fifo_full_140097941519888(0);
        
        fifo_inputs_140097941519944(0) <= outputs_140097941519888(0);
        outputs_full_140097941519888(0) <= fifo_full_140097941519944(0);
        
        fifo_inputs_140097941520000(0) <= outputs_140097941519944(0);
        outputs_full_140097941519944(0) <= fifo_full_140097941520000(0);
        
        fifo_inputs_140097941520056(0) <= outputs_140097941520000(0);
        outputs_full_140097941520000(0) <= fifo_full_140097941520056(0);
        
        fifo_inputs_140097941520112(0) <= outputs_140097941520056(0);
        outputs_full_140097941520056(0) <= fifo_full_140097941520112(0);
        
        fifo_inputs_140097941520168(0) <= outputs_140097941520112(0);
        outputs_full_140097941520112(0) <= fifo_full_140097941520168(0);
        
        fifo_inputs_140097941520224(0) <= outputs_140097941520168(0);
        outputs_full_140097941520168(0) <= fifo_full_140097941520224(0);
        
        fifo_inputs_140097941520280(0) <= outputs_140097941520224(0);
        outputs_full_140097941520224(0) <= fifo_full_140097941520280(0);
        
        fifo_inputs_140097941520336(0) <= outputs_140097941520280(0);
        outputs_full_140097941520280(0) <= fifo_full_140097941520336(0);
        
        fifo_inputs_140097941528648(0) <= outputs_140097941520336(0);
        outputs_full_140097941520336(0) <= fifo_full_140097941528648(0);
        
        fifo_inputs_140097941528704(0) <= outputs_140097941528648(0);
        outputs_full_140097941528648(0) <= fifo_full_140097941528704(0);
        
        fifo_inputs_140097941528760(0) <= outputs_140097941528704(0);
        outputs_full_140097941528704(0) <= fifo_full_140097941528760(0);
        
        fifo_inputs_140097941528816(0) <= outputs_140097941528760(0);
        outputs_full_140097941528760(0) <= fifo_full_140097941528816(0);
        
        fifo_inputs_140097941528872(0) <= outputs_140097941528816(0);
        outputs_full_140097941528816(0) <= fifo_full_140097941528872(0);
        
        fifo_inputs_140097941528928(0) <= outputs_140097941528872(0);
        outputs_full_140097941528872(0) <= fifo_full_140097941528928(0);
        
        fifo_inputs_140097941528984(0) <= outputs_140097941528928(0);
        outputs_full_140097941528928(0) <= fifo_full_140097941528984(0);
        
        fifo_inputs_140097941529040(0) <= outputs_140097941528984(0);
        outputs_full_140097941528984(0) <= fifo_full_140097941529040(0);
        
        fifo_inputs_140097941529096(0) <= outputs_140097941529040(0);
        outputs_full_140097941529040(0) <= fifo_full_140097941529096(0);
        
        fifo_inputs_140097941529152(0) <= outputs_140097941529096(0);
        outputs_full_140097941529096(0) <= fifo_full_140097941529152(0);
        
        fifo_inputs_140097941529208(0) <= outputs_140097941529152(0);
        outputs_full_140097941529152(0) <= fifo_full_140097941529208(0);
        
        fifo_inputs_140097941529264(0) <= outputs_140097941529208(0);
        outputs_full_140097941529208(0) <= fifo_full_140097941529264(0);
        
        fifo_inputs_140097941529320(0) <= outputs_140097941529264(0);
        outputs_full_140097941529264(0) <= fifo_full_140097941529320(0);
        
        fifo_inputs_140097941529376(0) <= outputs_140097941529320(0);
        outputs_full_140097941529320(0) <= fifo_full_140097941529376(0);
        
        fifo_inputs_140097941529432(0) <= outputs_140097941529376(0);
        outputs_full_140097941529376(0) <= fifo_full_140097941529432(0);
        
        fifo_inputs_140097941529488(0) <= outputs_140097941529432(0);
        outputs_full_140097941529432(0) <= fifo_full_140097941529488(0);
        
        fifo_inputs_140097941529544(0) <= outputs_140097941529488(0);
        outputs_full_140097941529488(0) <= fifo_full_140097941529544(0);
        
        fifo_inputs_140097941529600(0) <= outputs_140097941529544(0);
        outputs_full_140097941529544(0) <= fifo_full_140097941529600(0);
        
        fifo_inputs_140097941529656(0) <= outputs_140097941529600(0);
        outputs_full_140097941529600(0) <= fifo_full_140097941529656(0);
        
        fifo_inputs_140097941529712(0) <= outputs_140097941529656(0);
        outputs_full_140097941529656(0) <= fifo_full_140097941529712(0);
        
        fifo_inputs_140097941529768(0) <= outputs_140097941529712(0);
        outputs_full_140097941529712(0) <= fifo_full_140097941529768(0);
        
        fifo_inputs_140097941529824(0) <= outputs_140097941529768(0);
        outputs_full_140097941529768(0) <= fifo_full_140097941529824(0);
        
        fifo_inputs_140097941529880(0) <= outputs_140097941529824(0);
        outputs_full_140097941529824(0) <= fifo_full_140097941529880(0);
        
        fifo_inputs_140097941529936(0) <= outputs_140097941529880(0);
        outputs_full_140097941529880(0) <= fifo_full_140097941529936(0);
        
        fifo_inputs_140097941529992(0) <= outputs_140097941529936(0);
        outputs_full_140097941529936(0) <= fifo_full_140097941529992(0);
        
        fifo_inputs_140097941530048(0) <= outputs_140097941529992(0);
        outputs_full_140097941529992(0) <= fifo_full_140097941530048(0);
        
        fifo_inputs_140097941530104(0) <= outputs_140097941530048(0);
        outputs_full_140097941530048(0) <= fifo_full_140097941530104(0);
        
        fifo_inputs_140097941530160(0) <= outputs_140097941530104(0);
        outputs_full_140097941530104(0) <= fifo_full_140097941530160(0);
        
        fifo_inputs_140097941530216(0) <= outputs_140097941530160(0);
        outputs_full_140097941530160(0) <= fifo_full_140097941530216(0);
        
        fifo_inputs_140097941530272(0) <= outputs_140097941530216(0);
        outputs_full_140097941530216(0) <= fifo_full_140097941530272(0);
        
        fifo_inputs_140097941530328(0) <= outputs_140097941530272(0);
        outputs_full_140097941530272(0) <= fifo_full_140097941530328(0);
        
        fifo_inputs_140097941530384(0) <= outputs_140097941530328(0);
        outputs_full_140097941530328(0) <= fifo_full_140097941530384(0);
        
        fifo_inputs_140097941530440(0) <= outputs_140097941530384(0);
        outputs_full_140097941530384(0) <= fifo_full_140097941530440(0);
        
        fifo_inputs_140097941530496(0) <= outputs_140097941530440(0);
        outputs_full_140097941530440(0) <= fifo_full_140097941530496(0);
        
        fifo_inputs_140097941530552(0) <= outputs_140097941530496(0);
        outputs_full_140097941530496(0) <= fifo_full_140097941530552(0);
        
        fifo_inputs_140097941530608(0) <= outputs_140097941530552(0);
        outputs_full_140097941530552(0) <= fifo_full_140097941530608(0);
        
        fifo_inputs_140097941530664(0) <= outputs_140097941530608(0);
        outputs_full_140097941530608(0) <= fifo_full_140097941530664(0);
        
        fifo_inputs_140097941530720(0) <= outputs_140097941530664(0);
        outputs_full_140097941530664(0) <= fifo_full_140097941530720(0);
        
        fifo_inputs_140097941530776(0) <= outputs_140097941530720(0);
        outputs_full_140097941530720(0) <= fifo_full_140097941530776(0);
        
        fifo_inputs_140097941530832(0) <= outputs_140097941530776(0);
        outputs_full_140097941530776(0) <= fifo_full_140097941530832(0);
        
        fifo_inputs_140097941530888(0) <= outputs_140097941530832(0);
        outputs_full_140097941530832(0) <= fifo_full_140097941530888(0);
        
        fifo_inputs_140097941530944(0) <= outputs_140097941530888(0);
        outputs_full_140097941530888(0) <= fifo_full_140097941530944(0);
        
        fifo_inputs_140097941531000(0) <= outputs_140097941530944(0);
        outputs_full_140097941530944(0) <= fifo_full_140097941531000(0);
        
        fifo_inputs_140097941531056(0) <= outputs_140097941531000(0);
        outputs_full_140097941531000(0) <= fifo_full_140097941531056(0);
        
        fifo_inputs_140097941531112(0) <= outputs_140097941531056(0);
        outputs_full_140097941531056(0) <= fifo_full_140097941531112(0);
        
        fifo_inputs_140097941531168(0) <= outputs_140097941531112(0);
        outputs_full_140097941531112(0) <= fifo_full_140097941531168(0);
        
        fifo_inputs_140097941531224(0) <= outputs_140097941531168(0);
        outputs_full_140097941531168(0) <= fifo_full_140097941531224(0);
        
        fifo_inputs_140097941531280(0) <= outputs_140097941531224(0);
        outputs_full_140097941531224(0) <= fifo_full_140097941531280(0);
        
        fifo_inputs_140097941531336(0) <= outputs_140097941531280(0);
        outputs_full_140097941531280(0) <= fifo_full_140097941531336(0);
        
        fifo_inputs_140097941531392(0) <= outputs_140097941531336(0);
        outputs_full_140097941531336(0) <= fifo_full_140097941531392(0);
        
        fifo_inputs_140097941531448(0) <= outputs_140097941531392(0);
        outputs_full_140097941531392(0) <= fifo_full_140097941531448(0);
        
        fifo_inputs_140097941531504(0) <= outputs_140097941531448(0);
        outputs_full_140097941531448(0) <= fifo_full_140097941531504(0);
        
        fifo_inputs_140097941531560(0) <= outputs_140097941531504(0);
        outputs_full_140097941531504(0) <= fifo_full_140097941531560(0);
        
        fifo_inputs_140097941531616(0) <= outputs_140097941531560(0);
        outputs_full_140097941531560(0) <= fifo_full_140097941531616(0);
        
        fifo_inputs_140097941531672(0) <= outputs_140097941531616(0);
        outputs_full_140097941531616(0) <= fifo_full_140097941531672(0);
        
        fifo_inputs_140097941531728(0) <= outputs_140097941531672(0);
        outputs_full_140097941531672(0) <= fifo_full_140097941531728(0);
        
        fifo_inputs_140097941531784(0) <= outputs_140097941531728(0);
        outputs_full_140097941531728(0) <= fifo_full_140097941531784(0);
        
        fifo_inputs_140097941531840(0) <= outputs_140097941531784(0);
        outputs_full_140097941531784(0) <= fifo_full_140097941531840(0);
        
        fifo_inputs_140097941531896(0) <= outputs_140097941531840(0);
        outputs_full_140097941531840(0) <= fifo_full_140097941531896(0);
        
        fifo_inputs_140097941531952(0) <= outputs_140097941531896(0);
        outputs_full_140097941531896(0) <= fifo_full_140097941531952(0);
        
        fifo_inputs_140097941532008(0) <= outputs_140097941531952(0);
        outputs_full_140097941531952(0) <= fifo_full_140097941532008(0);
        
        fifo_inputs_140097941532064(0) <= outputs_140097941532008(0);
        outputs_full_140097941532008(0) <= fifo_full_140097941532064(0);
        
        fifo_inputs_140097941532120(0) <= outputs_140097941532064(0);
        outputs_full_140097941532064(0) <= fifo_full_140097941532120(0);
        
        fifo_inputs_140097941532176(0) <= outputs_140097941532120(0);
        outputs_full_140097941532120(0) <= fifo_full_140097941532176(0);
        
        fifo_inputs_140097941532232(0) <= outputs_140097941532176(0);
        outputs_full_140097941532176(0) <= fifo_full_140097941532232(0);
        
        fifo_inputs_140097941532288(0) <= outputs_140097941532232(0);
        outputs_full_140097941532232(0) <= fifo_full_140097941532288(0);
        
        fifo_inputs_140097941532344(0) <= outputs_140097941532288(0);
        outputs_full_140097941532288(0) <= fifo_full_140097941532344(0);
        
        fifo_inputs_140097941532400(0) <= outputs_140097941532344(0);
        outputs_full_140097941532344(0) <= fifo_full_140097941532400(0);
        
        fifo_inputs_140097941532456(0) <= outputs_140097941532400(0);
        outputs_full_140097941532400(0) <= fifo_full_140097941532456(0);
        
        fifo_inputs_140097941532512(0) <= outputs_140097941532456(0);
        outputs_full_140097941532456(0) <= fifo_full_140097941532512(0);
        
        fifo_inputs_140097941532568(0) <= outputs_140097941532512(0);
        outputs_full_140097941532512(0) <= fifo_full_140097941532568(0);
        
        fifo_inputs_140097941532624(0) <= outputs_140097941532568(0);
        outputs_full_140097941532568(0) <= fifo_full_140097941532624(0);
        
        fifo_inputs_140097941540936(0) <= outputs_140097941532624(0);
        outputs_full_140097941532624(0) <= fifo_full_140097941540936(0);
        
        fifo_inputs_140097941540992(0) <= outputs_140097941540936(0);
        outputs_full_140097941540936(0) <= fifo_full_140097941540992(0);
        
        fifo_inputs_140097941541048(0) <= outputs_140097941540992(0);
        outputs_full_140097941540992(0) <= fifo_full_140097941541048(0);
        
        fifo_inputs_140097941541104(0) <= outputs_140097941541048(0);
        outputs_full_140097941541048(0) <= fifo_full_140097941541104(0);
        
        fifo_inputs_140097941541160(0) <= outputs_140097941541104(0);
        outputs_full_140097941541104(0) <= fifo_full_140097941541160(0);
        
        fifo_inputs_140097941541216(0) <= outputs_140097941541160(0);
        outputs_full_140097941541160(0) <= fifo_full_140097941541216(0);
        
        fifo_inputs_140097941541272(0) <= outputs_140097941541216(0);
        outputs_full_140097941541216(0) <= fifo_full_140097941541272(0);
        
        fifo_inputs_140097941541328(0) <= outputs_140097941541272(0);
        outputs_full_140097941541272(0) <= fifo_full_140097941541328(0);
        
        fifo_inputs_140097941541384(0) <= outputs_140097941541328(0);
        outputs_full_140097941541328(0) <= fifo_full_140097941541384(0);
        
        fifo_inputs_140097941541440(0) <= outputs_140097941541384(0);
        outputs_full_140097941541384(0) <= fifo_full_140097941541440(0);
        
        fifo_inputs_140097941541496(0) <= outputs_140097941541440(0);
        outputs_full_140097941541440(0) <= fifo_full_140097941541496(0);
        
        fifo_inputs_140097941541552(0) <= outputs_140097941541496(0);
        outputs_full_140097941541496(0) <= fifo_full_140097941541552(0);
        
        fifo_inputs_140097941541608(0) <= outputs_140097941541552(0);
        outputs_full_140097941541552(0) <= fifo_full_140097941541608(0);
        
        fifo_inputs_140097941541664(0) <= outputs_140097941541608(0);
        outputs_full_140097941541608(0) <= fifo_full_140097941541664(0);
        
        fifo_inputs_140097941541720(0) <= outputs_140097941541664(0);
        outputs_full_140097941541664(0) <= fifo_full_140097941541720(0);
        
        fifo_inputs_140097941541776(0) <= outputs_140097941541720(0);
        outputs_full_140097941541720(0) <= fifo_full_140097941541776(0);
        
        fifo_inputs_140097941541832(0) <= outputs_140097941541776(0);
        outputs_full_140097941541776(0) <= fifo_full_140097941541832(0);
        
        fifo_inputs_140097941541888(0) <= outputs_140097941541832(0);
        outputs_full_140097941541832(0) <= fifo_full_140097941541888(0);
        
        fifo_inputs_140097941541944(0) <= outputs_140097941541888(0);
        outputs_full_140097941541888(0) <= fifo_full_140097941541944(0);
        
        fifo_inputs_140097941542000(0) <= outputs_140097941541944(0);
        outputs_full_140097941541944(0) <= fifo_full_140097941542000(0);
        
        fifo_inputs_140097941542056(0) <= outputs_140097941542000(0);
        outputs_full_140097941542000(0) <= fifo_full_140097941542056(0);
        
        fifo_inputs_140097941542112(0) <= outputs_140097941542056(0);
        outputs_full_140097941542056(0) <= fifo_full_140097941542112(0);
        
        fifo_inputs_140097941542168(0) <= outputs_140097941542112(0);
        outputs_full_140097941542112(0) <= fifo_full_140097941542168(0);
        
        fifo_inputs_140097941542224(0) <= outputs_140097941542168(0);
        outputs_full_140097941542168(0) <= fifo_full_140097941542224(0);
        
        fifo_inputs_140097941542280(0) <= outputs_140097941542224(0);
        outputs_full_140097941542224(0) <= fifo_full_140097941542280(0);
        
        fifo_inputs_140097941542336(0) <= outputs_140097941542280(0);
        outputs_full_140097941542280(0) <= fifo_full_140097941542336(0);
        
        fifo_inputs_140097941542392(0) <= outputs_140097941542336(0);
        outputs_full_140097941542336(0) <= fifo_full_140097941542392(0);
        
        fifo_inputs_140097941542448(0) <= outputs_140097941542392(0);
        outputs_full_140097941542392(0) <= fifo_full_140097941542448(0);
        
        fifo_inputs_140097941542504(0) <= outputs_140097941542448(0);
        outputs_full_140097941542448(0) <= fifo_full_140097941542504(0);
        
        fifo_inputs_140097941542560(0) <= outputs_140097941542504(0);
        outputs_full_140097941542504(0) <= fifo_full_140097941542560(0);
        
        fifo_inputs_140097941542616(0) <= outputs_140097941542560(0);
        outputs_full_140097941542560(0) <= fifo_full_140097941542616(0);
        
        fifo_inputs_140097941542672(0) <= outputs_140097941542616(0);
        outputs_full_140097941542616(0) <= fifo_full_140097941542672(0);
        
        fifo_inputs_140097941542728(0) <= outputs_140097941542672(0);
        outputs_full_140097941542672(0) <= fifo_full_140097941542728(0);
        
        fifo_inputs_140097941542784(0) <= outputs_140097941542728(0);
        outputs_full_140097941542728(0) <= fifo_full_140097941542784(0);
        
        fifo_inputs_140097941542840(0) <= outputs_140097941542784(0);
        outputs_full_140097941542784(0) <= fifo_full_140097941542840(0);
        
        fifo_inputs_140097941542896(0) <= outputs_140097941542840(0);
        outputs_full_140097941542840(0) <= fifo_full_140097941542896(0);
        
        fifo_inputs_140097941542952(0) <= outputs_140097941542896(0);
        outputs_full_140097941542896(0) <= fifo_full_140097941542952(0);
        
        fifo_inputs_140097941543008(0) <= outputs_140097941542952(0);
        outputs_full_140097941542952(0) <= fifo_full_140097941543008(0);
        
        fifo_inputs_140097941543064(0) <= outputs_140097941543008(0);
        outputs_full_140097941543008(0) <= fifo_full_140097941543064(0);
        
        fifo_inputs_140097941543120(0) <= outputs_140097941543064(0);
        outputs_full_140097941543064(0) <= fifo_full_140097941543120(0);
        
        fifo_inputs_140097941543176(0) <= outputs_140097941543120(0);
        outputs_full_140097941543120(0) <= fifo_full_140097941543176(0);
        
        fifo_inputs_140097941543232(0) <= outputs_140097941543176(0);
        outputs_full_140097941543176(0) <= fifo_full_140097941543232(0);
        
        fifo_inputs_140097941543288(0) <= outputs_140097941543232(0);
        outputs_full_140097941543232(0) <= fifo_full_140097941543288(0);
        
        fifo_inputs_140097941543344(0) <= outputs_140097941543288(0);
        outputs_full_140097941543288(0) <= fifo_full_140097941543344(0);
        
        fifo_inputs_140097941543400(0) <= outputs_140097941543344(0);
        outputs_full_140097941543344(0) <= fifo_full_140097941543400(0);
        
        fifo_inputs_140097941543456(0) <= outputs_140097941543400(0);
        outputs_full_140097941543400(0) <= fifo_full_140097941543456(0);
        
        fifo_inputs_140097941543512(0) <= outputs_140097941543456(0);
        outputs_full_140097941543456(0) <= fifo_full_140097941543512(0);
        
        fifo_inputs_140097941543568(0) <= outputs_140097941543512(0);
        outputs_full_140097941543512(0) <= fifo_full_140097941543568(0);
        
        fifo_inputs_140097941543624(0) <= outputs_140097941543568(0);
        outputs_full_140097941543568(0) <= fifo_full_140097941543624(0);
        
        fifo_inputs_140097941543680(0) <= outputs_140097941543624(0);
        outputs_full_140097941543624(0) <= fifo_full_140097941543680(0);
        
        fifo_inputs_140097941543736(0) <= outputs_140097941543680(0);
        outputs_full_140097941543680(0) <= fifo_full_140097941543736(0);
        
        fifo_inputs_140097941543792(0) <= outputs_140097941543736(0);
        outputs_full_140097941543736(0) <= fifo_full_140097941543792(0);
        
        fifo_inputs_140097941543848(0) <= outputs_140097941543792(0);
        outputs_full_140097941543792(0) <= fifo_full_140097941543848(0);
        
        fifo_inputs_140097941543904(0) <= outputs_140097941543848(0);
        outputs_full_140097941543848(0) <= fifo_full_140097941543904(0);
        
        fifo_inputs_140097941543960(0) <= outputs_140097941543904(0);
        outputs_full_140097941543904(0) <= fifo_full_140097941543960(0);
        
        fifo_inputs_140097941544016(0) <= outputs_140097941543960(0);
        outputs_full_140097941543960(0) <= fifo_full_140097941544016(0);
        
        fifo_inputs_140097941544072(0) <= outputs_140097941544016(0);
        outputs_full_140097941544016(0) <= fifo_full_140097941544072(0);
        
        fifo_inputs_140097941544128(0) <= outputs_140097941544072(0);
        outputs_full_140097941544072(0) <= fifo_full_140097941544128(0);
        
        fifo_inputs_140097941544184(0) <= outputs_140097941544128(0);
        outputs_full_140097941544128(0) <= fifo_full_140097941544184(0);
        
        fifo_inputs_140097941544240(0) <= outputs_140097941544184(0);
        outputs_full_140097941544184(0) <= fifo_full_140097941544240(0);
        
        fifo_inputs_140097941544296(0) <= outputs_140097941544240(0);
        outputs_full_140097941544240(0) <= fifo_full_140097941544296(0);
        
        fifo_inputs_140097941544352(0) <= outputs_140097941544296(0);
        outputs_full_140097941544296(0) <= fifo_full_140097941544352(0);
        
        fifo_inputs_140097941544408(0) <= outputs_140097941544352(0);
        outputs_full_140097941544352(0) <= fifo_full_140097941544408(0);
        
        fifo_inputs_140097941544464(0) <= outputs_140097941544408(0);
        outputs_full_140097941544408(0) <= fifo_full_140097941544464(0);
        
        fifo_inputs_140097941544520(0) <= outputs_140097941544464(0);
        outputs_full_140097941544464(0) <= fifo_full_140097941544520(0);
        
        fifo_inputs_140097941544576(0) <= outputs_140097941544520(0);
        outputs_full_140097941544520(0) <= fifo_full_140097941544576(0);
        
        fifo_inputs_140097941544632(0) <= outputs_140097941544576(0);
        outputs_full_140097941544576(0) <= fifo_full_140097941544632(0);
        
        fifo_inputs_140097941544688(0) <= outputs_140097941544632(0);
        outputs_full_140097941544632(0) <= fifo_full_140097941544688(0);
        
        fifo_inputs_140097941544744(0) <= outputs_140097941544688(0);
        outputs_full_140097941544688(0) <= fifo_full_140097941544744(0);
        
        fifo_inputs_140097941544800(0) <= outputs_140097941544744(0);
        outputs_full_140097941544744(0) <= fifo_full_140097941544800(0);
        
        fifo_inputs_140097941544856(0) <= outputs_140097941544800(0);
        outputs_full_140097941544800(0) <= fifo_full_140097941544856(0);
        
        fifo_inputs_140097941544912(0) <= outputs_140097941544856(0);
        outputs_full_140097941544856(0) <= fifo_full_140097941544912(0);
        
        fifo_inputs_140097941553224(0) <= outputs_140097941544912(0);
        outputs_full_140097941544912(0) <= fifo_full_140097941553224(0);
        
        fifo_inputs_140097941553280(0) <= outputs_140097941553224(0);
        outputs_full_140097941553224(0) <= fifo_full_140097941553280(0);
        
        fifo_inputs_140097941553336(0) <= outputs_140097941553280(0);
        outputs_full_140097941553280(0) <= fifo_full_140097941553336(0);
        
        fifo_inputs_140097941553392(0) <= outputs_140097941553336(0);
        outputs_full_140097941553336(0) <= fifo_full_140097941553392(0);
        
        fifo_inputs_140097941553448(0) <= outputs_140097941553392(0);
        outputs_full_140097941553392(0) <= fifo_full_140097941553448(0);
        
        fifo_inputs_140097941553504(0) <= outputs_140097941553448(0);
        outputs_full_140097941553448(0) <= fifo_full_140097941553504(0);
        
        fifo_inputs_140097941553560(0) <= outputs_140097941553504(0);
        outputs_full_140097941553504(0) <= fifo_full_140097941553560(0);
        
        fifo_inputs_140097941553616(0) <= outputs_140097941553560(0);
        outputs_full_140097941553560(0) <= fifo_full_140097941553616(0);
        
        fifo_inputs_140097941553672(0) <= outputs_140097941553616(0);
        outputs_full_140097941553616(0) <= fifo_full_140097941553672(0);
        
        fifo_inputs_140097941553728(0) <= outputs_140097941553672(0);
        outputs_full_140097941553672(0) <= fifo_full_140097941553728(0);
        
        fifo_inputs_140097941553784(0) <= outputs_140097941553728(0);
        outputs_full_140097941553728(0) <= fifo_full_140097941553784(0);
        
        fifo_inputs_140097941553840(0) <= outputs_140097941553784(0);
        outputs_full_140097941553784(0) <= fifo_full_140097941553840(0);
        
        fifo_inputs_140097941553896(0) <= outputs_140097941553840(0);
        outputs_full_140097941553840(0) <= fifo_full_140097941553896(0);
        
        fifo_inputs_140097941553952(0) <= outputs_140097941553896(0);
        outputs_full_140097941553896(0) <= fifo_full_140097941553952(0);
        
        fifo_inputs_140097941554008(0) <= outputs_140097941553952(0);
        outputs_full_140097941553952(0) <= fifo_full_140097941554008(0);
        
        fifo_inputs_140097941554064(0) <= outputs_140097941554008(0);
        outputs_full_140097941554008(0) <= fifo_full_140097941554064(0);
        
        fifo_inputs_140097941554120(0) <= outputs_140097941554064(0);
        outputs_full_140097941554064(0) <= fifo_full_140097941554120(0);
        
        fifo_inputs_140097941554176(0) <= outputs_140097941554120(0);
        outputs_full_140097941554120(0) <= fifo_full_140097941554176(0);
        
        fifo_inputs_140097941554232(0) <= outputs_140097941554176(0);
        outputs_full_140097941554176(0) <= fifo_full_140097941554232(0);
        
        fifo_inputs_140097941554288(0) <= outputs_140097941554232(0);
        outputs_full_140097941554232(0) <= fifo_full_140097941554288(0);
        
        fifo_inputs_140097941554344(0) <= outputs_140097941554288(0);
        outputs_full_140097941554288(0) <= fifo_full_140097941554344(0);
        
        fifo_inputs_140097941554400(0) <= outputs_140097941554344(0);
        outputs_full_140097941554344(0) <= fifo_full_140097941554400(0);
        
        fifo_inputs_140097941554456(0) <= outputs_140097941554400(0);
        outputs_full_140097941554400(0) <= fifo_full_140097941554456(0);
        
        fifo_inputs_140097941554512(0) <= outputs_140097941554456(0);
        outputs_full_140097941554456(0) <= fifo_full_140097941554512(0);
        
        fifo_inputs_140097941554568(0) <= outputs_140097941554512(0);
        outputs_full_140097941554512(0) <= fifo_full_140097941554568(0);
        
        fifo_inputs_140097941554624(0) <= outputs_140097941554568(0);
        outputs_full_140097941554568(0) <= fifo_full_140097941554624(0);
        
        fifo_inputs_140097941554680(0) <= outputs_140097941554624(0);
        outputs_full_140097941554624(0) <= fifo_full_140097941554680(0);
        
        fifo_inputs_140097941554736(0) <= outputs_140097941554680(0);
        outputs_full_140097941554680(0) <= fifo_full_140097941554736(0);
        
        fifo_inputs_140097941554792(0) <= outputs_140097941554736(0);
        outputs_full_140097941554736(0) <= fifo_full_140097941554792(0);
        
        fifo_inputs_140097941554848(0) <= outputs_140097941554792(0);
        outputs_full_140097941554792(0) <= fifo_full_140097941554848(0);
        
        fifo_inputs_140097941554904(0) <= outputs_140097941554848(0);
        outputs_full_140097941554848(0) <= fifo_full_140097941554904(0);
        
        fifo_inputs_140097941554960(0) <= outputs_140097941554904(0);
        outputs_full_140097941554904(0) <= fifo_full_140097941554960(0);
        
        fifo_inputs_140097941555016(0) <= outputs_140097941554960(0);
        outputs_full_140097941554960(0) <= fifo_full_140097941555016(0);
        
        fifo_inputs_140097941555072(0) <= outputs_140097941555016(0);
        outputs_full_140097941555016(0) <= fifo_full_140097941555072(0);
        
        fifo_inputs_140097941555128(0) <= outputs_140097941555072(0);
        outputs_full_140097941555072(0) <= fifo_full_140097941555128(0);
        
        fifo_inputs_140097941555184(0) <= outputs_140097941555128(0);
        outputs_full_140097941555128(0) <= fifo_full_140097941555184(0);
        
        fifo_inputs_140097941555240(0) <= outputs_140097941555184(0);
        outputs_full_140097941555184(0) <= fifo_full_140097941555240(0);
        
        fifo_inputs_140097941555296(0) <= outputs_140097941555240(0);
        outputs_full_140097941555240(0) <= fifo_full_140097941555296(0);
        
        fifo_inputs_140097941555352(0) <= outputs_140097941555296(0);
        outputs_full_140097941555296(0) <= fifo_full_140097941555352(0);
        
        fifo_inputs_140097941555408(0) <= outputs_140097941555352(0);
        outputs_full_140097941555352(0) <= fifo_full_140097941555408(0);
        
        fifo_inputs_140097941555464(0) <= outputs_140097941555408(0);
        outputs_full_140097941555408(0) <= fifo_full_140097941555464(0);
        
        fifo_inputs_140097941555520(0) <= outputs_140097941555464(0);
        outputs_full_140097941555464(0) <= fifo_full_140097941555520(0);
        
        fifo_inputs_140097941555576(0) <= outputs_140097941555520(0);
        outputs_full_140097941555520(0) <= fifo_full_140097941555576(0);
        
        fifo_inputs_140097941555632(0) <= outputs_140097941555576(0);
        outputs_full_140097941555576(0) <= fifo_full_140097941555632(0);
        
        fifo_inputs_140097941555688(0) <= outputs_140097941555632(0);
        outputs_full_140097941555632(0) <= fifo_full_140097941555688(0);
        

    
        core_inst_140097944041960: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944041960,
            fifo_full => fifo_full_140097944041960,
            outputs => outputs_140097944041960,
            outputs_full => outputs_full_140097944041960
        );
        
        core_inst_140097944041904: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944041904,
            fifo_full => fifo_full_140097944041904,
            outputs => outputs_140097944041904,
            outputs_full => outputs_full_140097944041904
        );
        
        core_inst_140097944042128: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944042128,
            fifo_full => fifo_full_140097944042128,
            outputs => outputs_140097944042128,
            outputs_full => outputs_full_140097944042128
        );
        
        core_inst_140097944042072: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944042072,
            fifo_full => fifo_full_140097944042072,
            outputs => outputs_140097944042072,
            outputs_full => outputs_full_140097944042072
        );
        
        core_inst_140097944042184: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944042184,
            fifo_full => fifo_full_140097944042184,
            outputs => outputs_140097944042184,
            outputs_full => outputs_full_140097944042184
        );
        
        core_inst_140097944042240: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944042240,
            fifo_full => fifo_full_140097944042240,
            outputs => outputs_140097944042240,
            outputs_full => outputs_full_140097944042240
        );
        
        core_inst_140097944042296: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944042296,
            fifo_full => fifo_full_140097944042296,
            outputs => outputs_140097944042296,
            outputs_full => outputs_full_140097944042296
        );
        
        core_inst_140097944042352: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944042352,
            fifo_full => fifo_full_140097944042352,
            outputs => outputs_140097944042352,
            outputs_full => outputs_full_140097944042352
        );
        
        core_inst_140097944042408: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944042408,
            fifo_full => fifo_full_140097944042408,
            outputs => outputs_140097944042408,
            outputs_full => outputs_full_140097944042408
        );
        
        core_inst_140097944042464: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944042464,
            fifo_full => fifo_full_140097944042464,
            outputs => outputs_140097944042464,
            outputs_full => outputs_full_140097944042464
        );
        
        core_inst_140097944042016: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944042016,
            fifo_full => fifo_full_140097944042016,
            outputs => outputs_140097944042016,
            outputs_full => outputs_full_140097944042016
        );
        
        core_inst_140097944042520: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944042520,
            fifo_full => fifo_full_140097944042520,
            outputs => outputs_140097944042520,
            outputs_full => outputs_full_140097944042520
        );
        
        core_inst_140097944042576: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944042576,
            fifo_full => fifo_full_140097944042576,
            outputs => outputs_140097944042576,
            outputs_full => outputs_full_140097944042576
        );
        
        core_inst_140097944042632: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944042632,
            fifo_full => fifo_full_140097944042632,
            outputs => outputs_140097944042632,
            outputs_full => outputs_full_140097944042632
        );
        
        core_inst_140097944042688: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944042688,
            fifo_full => fifo_full_140097944042688,
            outputs => outputs_140097944042688,
            outputs_full => outputs_full_140097944042688
        );
        
        core_inst_140097944042744: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944042744,
            fifo_full => fifo_full_140097944042744,
            outputs => outputs_140097944042744,
            outputs_full => outputs_full_140097944042744
        );
        
        core_inst_140097944042800: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944042800,
            fifo_full => fifo_full_140097944042800,
            outputs => outputs_140097944042800,
            outputs_full => outputs_full_140097944042800
        );
        
        core_inst_140097944042856: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944042856,
            fifo_full => fifo_full_140097944042856,
            outputs => outputs_140097944042856,
            outputs_full => outputs_full_140097944042856
        );
        
        core_inst_140097944042912: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944042912,
            fifo_full => fifo_full_140097944042912,
            outputs => outputs_140097944042912,
            outputs_full => outputs_full_140097944042912
        );
        
        core_inst_140097944042968: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944042968,
            fifo_full => fifo_full_140097944042968,
            outputs => outputs_140097944042968,
            outputs_full => outputs_full_140097944042968
        );
        
        core_inst_140097944043024: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944043024,
            fifo_full => fifo_full_140097944043024,
            outputs => outputs_140097944043024,
            outputs_full => outputs_full_140097944043024
        );
        
        core_inst_140097944043080: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944043080,
            fifo_full => fifo_full_140097944043080,
            outputs => outputs_140097944043080,
            outputs_full => outputs_full_140097944043080
        );
        
        core_inst_140097944043136: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944043136,
            fifo_full => fifo_full_140097944043136,
            outputs => outputs_140097944043136,
            outputs_full => outputs_full_140097944043136
        );
        
        core_inst_140097944043192: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944043192,
            fifo_full => fifo_full_140097944043192,
            outputs => outputs_140097944043192,
            outputs_full => outputs_full_140097944043192
        );
        
        core_inst_140097944043248: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944043248,
            fifo_full => fifo_full_140097944043248,
            outputs => outputs_140097944043248,
            outputs_full => outputs_full_140097944043248
        );
        
        core_inst_140097944043304: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944043304,
            fifo_full => fifo_full_140097944043304,
            outputs => outputs_140097944043304,
            outputs_full => outputs_full_140097944043304
        );
        
        core_inst_140097944043360: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944043360,
            fifo_full => fifo_full_140097944043360,
            outputs => outputs_140097944043360,
            outputs_full => outputs_full_140097944043360
        );
        
        core_inst_140097944043416: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944043416,
            fifo_full => fifo_full_140097944043416,
            outputs => outputs_140097944043416,
            outputs_full => outputs_full_140097944043416
        );
        
        core_inst_140097944043472: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944043472,
            fifo_full => fifo_full_140097944043472,
            outputs => outputs_140097944043472,
            outputs_full => outputs_full_140097944043472
        );
        
        core_inst_140097944076360: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944076360,
            fifo_full => fifo_full_140097944076360,
            outputs => outputs_140097944076360,
            outputs_full => outputs_full_140097944076360
        );
        
        core_inst_140097944076416: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944076416,
            fifo_full => fifo_full_140097944076416,
            outputs => outputs_140097944076416,
            outputs_full => outputs_full_140097944076416
        );
        
        core_inst_140097944076472: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944076472,
            fifo_full => fifo_full_140097944076472,
            outputs => outputs_140097944076472,
            outputs_full => outputs_full_140097944076472
        );
        
        core_inst_140097944076528: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944076528,
            fifo_full => fifo_full_140097944076528,
            outputs => outputs_140097944076528,
            outputs_full => outputs_full_140097944076528
        );
        
        core_inst_140097944076584: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944076584,
            fifo_full => fifo_full_140097944076584,
            outputs => outputs_140097944076584,
            outputs_full => outputs_full_140097944076584
        );
        
        core_inst_140097944076640: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944076640,
            fifo_full => fifo_full_140097944076640,
            outputs => outputs_140097944076640,
            outputs_full => outputs_full_140097944076640
        );
        
        core_inst_140097944076696: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944076696,
            fifo_full => fifo_full_140097944076696,
            outputs => outputs_140097944076696,
            outputs_full => outputs_full_140097944076696
        );
        
        core_inst_140097944076752: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944076752,
            fifo_full => fifo_full_140097944076752,
            outputs => outputs_140097944076752,
            outputs_full => outputs_full_140097944076752
        );
        
        core_inst_140097944076808: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944076808,
            fifo_full => fifo_full_140097944076808,
            outputs => outputs_140097944076808,
            outputs_full => outputs_full_140097944076808
        );
        
        core_inst_140097944076864: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944076864,
            fifo_full => fifo_full_140097944076864,
            outputs => outputs_140097944076864,
            outputs_full => outputs_full_140097944076864
        );
        
        core_inst_140097944076920: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944076920,
            fifo_full => fifo_full_140097944076920,
            outputs => outputs_140097944076920,
            outputs_full => outputs_full_140097944076920
        );
        
        core_inst_140097944076976: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944076976,
            fifo_full => fifo_full_140097944076976,
            outputs => outputs_140097944076976,
            outputs_full => outputs_full_140097944076976
        );
        
        core_inst_140097944077032: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944077032,
            fifo_full => fifo_full_140097944077032,
            outputs => outputs_140097944077032,
            outputs_full => outputs_full_140097944077032
        );
        
        core_inst_140097944077088: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944077088,
            fifo_full => fifo_full_140097944077088,
            outputs => outputs_140097944077088,
            outputs_full => outputs_full_140097944077088
        );
        
        core_inst_140097944077144: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944077144,
            fifo_full => fifo_full_140097944077144,
            outputs => outputs_140097944077144,
            outputs_full => outputs_full_140097944077144
        );
        
        core_inst_140097944077200: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944077200,
            fifo_full => fifo_full_140097944077200,
            outputs => outputs_140097944077200,
            outputs_full => outputs_full_140097944077200
        );
        
        core_inst_140097944077256: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944077256,
            fifo_full => fifo_full_140097944077256,
            outputs => outputs_140097944077256,
            outputs_full => outputs_full_140097944077256
        );
        
        core_inst_140097944077312: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944077312,
            fifo_full => fifo_full_140097944077312,
            outputs => outputs_140097944077312,
            outputs_full => outputs_full_140097944077312
        );
        
        core_inst_140097944077368: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944077368,
            fifo_full => fifo_full_140097944077368,
            outputs => outputs_140097944077368,
            outputs_full => outputs_full_140097944077368
        );
        
        core_inst_140097944077424: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944077424,
            fifo_full => fifo_full_140097944077424,
            outputs => outputs_140097944077424,
            outputs_full => outputs_full_140097944077424
        );
        
        core_inst_140097944077480: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944077480,
            fifo_full => fifo_full_140097944077480,
            outputs => outputs_140097944077480,
            outputs_full => outputs_full_140097944077480
        );
        
        core_inst_140097944077536: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944077536,
            fifo_full => fifo_full_140097944077536,
            outputs => outputs_140097944077536,
            outputs_full => outputs_full_140097944077536
        );
        
        core_inst_140097944077592: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944077592,
            fifo_full => fifo_full_140097944077592,
            outputs => outputs_140097944077592,
            outputs_full => outputs_full_140097944077592
        );
        
        core_inst_140097944077648: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944077648,
            fifo_full => fifo_full_140097944077648,
            outputs => outputs_140097944077648,
            outputs_full => outputs_full_140097944077648
        );
        
        core_inst_140097944077704: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944077704,
            fifo_full => fifo_full_140097944077704,
            outputs => outputs_140097944077704,
            outputs_full => outputs_full_140097944077704
        );
        
        core_inst_140097944077760: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944077760,
            fifo_full => fifo_full_140097944077760,
            outputs => outputs_140097944077760,
            outputs_full => outputs_full_140097944077760
        );
        
        core_inst_140097944077816: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944077816,
            fifo_full => fifo_full_140097944077816,
            outputs => outputs_140097944077816,
            outputs_full => outputs_full_140097944077816
        );
        
        core_inst_140097944077872: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944077872,
            fifo_full => fifo_full_140097944077872,
            outputs => outputs_140097944077872,
            outputs_full => outputs_full_140097944077872
        );
        
        core_inst_140097944077928: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944077928,
            fifo_full => fifo_full_140097944077928,
            outputs => outputs_140097944077928,
            outputs_full => outputs_full_140097944077928
        );
        
        core_inst_140097944077984: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944077984,
            fifo_full => fifo_full_140097944077984,
            outputs => outputs_140097944077984,
            outputs_full => outputs_full_140097944077984
        );
        
        core_inst_140097944078040: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944078040,
            fifo_full => fifo_full_140097944078040,
            outputs => outputs_140097944078040,
            outputs_full => outputs_full_140097944078040
        );
        
        core_inst_140097944078096: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944078096,
            fifo_full => fifo_full_140097944078096,
            outputs => outputs_140097944078096,
            outputs_full => outputs_full_140097944078096
        );
        
        core_inst_140097944078152: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944078152,
            fifo_full => fifo_full_140097944078152,
            outputs => outputs_140097944078152,
            outputs_full => outputs_full_140097944078152
        );
        
        core_inst_140097944078208: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944078208,
            fifo_full => fifo_full_140097944078208,
            outputs => outputs_140097944078208,
            outputs_full => outputs_full_140097944078208
        );
        
        core_inst_140097944078264: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944078264,
            fifo_full => fifo_full_140097944078264,
            outputs => outputs_140097944078264,
            outputs_full => outputs_full_140097944078264
        );
        
        core_inst_140097944078320: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944078320,
            fifo_full => fifo_full_140097944078320,
            outputs => outputs_140097944078320,
            outputs_full => outputs_full_140097944078320
        );
        
        core_inst_140097944078376: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944078376,
            fifo_full => fifo_full_140097944078376,
            outputs => outputs_140097944078376,
            outputs_full => outputs_full_140097944078376
        );
        
        core_inst_140097944078432: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944078432,
            fifo_full => fifo_full_140097944078432,
            outputs => outputs_140097944078432,
            outputs_full => outputs_full_140097944078432
        );
        
        core_inst_140097944078488: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944078488,
            fifo_full => fifo_full_140097944078488,
            outputs => outputs_140097944078488,
            outputs_full => outputs_full_140097944078488
        );
        
        core_inst_140097944078544: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944078544,
            fifo_full => fifo_full_140097944078544,
            outputs => outputs_140097944078544,
            outputs_full => outputs_full_140097944078544
        );
        
        core_inst_140097944078600: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944078600,
            fifo_full => fifo_full_140097944078600,
            outputs => outputs_140097944078600,
            outputs_full => outputs_full_140097944078600
        );
        
        core_inst_140097944078656: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944078656,
            fifo_full => fifo_full_140097944078656,
            outputs => outputs_140097944078656,
            outputs_full => outputs_full_140097944078656
        );
        
        core_inst_140097944078712: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944078712,
            fifo_full => fifo_full_140097944078712,
            outputs => outputs_140097944078712,
            outputs_full => outputs_full_140097944078712
        );
        
        core_inst_140097944078768: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944078768,
            fifo_full => fifo_full_140097944078768,
            outputs => outputs_140097944078768,
            outputs_full => outputs_full_140097944078768
        );
        
        core_inst_140097944078824: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944078824,
            fifo_full => fifo_full_140097944078824,
            outputs => outputs_140097944078824,
            outputs_full => outputs_full_140097944078824
        );
        
        core_inst_140097944078880: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944078880,
            fifo_full => fifo_full_140097944078880,
            outputs => outputs_140097944078880,
            outputs_full => outputs_full_140097944078880
        );
        
        core_inst_140097944078936: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944078936,
            fifo_full => fifo_full_140097944078936,
            outputs => outputs_140097944078936,
            outputs_full => outputs_full_140097944078936
        );
        
        core_inst_140097944078992: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944078992,
            fifo_full => fifo_full_140097944078992,
            outputs => outputs_140097944078992,
            outputs_full => outputs_full_140097944078992
        );
        
        core_inst_140097944079048: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944079048,
            fifo_full => fifo_full_140097944079048,
            outputs => outputs_140097944079048,
            outputs_full => outputs_full_140097944079048
        );
        
        core_inst_140097944079104: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944079104,
            fifo_full => fifo_full_140097944079104,
            outputs => outputs_140097944079104,
            outputs_full => outputs_full_140097944079104
        );
        
        core_inst_140097944079160: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944079160,
            fifo_full => fifo_full_140097944079160,
            outputs => outputs_140097944079160,
            outputs_full => outputs_full_140097944079160
        );
        
        core_inst_140097944079216: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944079216,
            fifo_full => fifo_full_140097944079216,
            outputs => outputs_140097944079216,
            outputs_full => outputs_full_140097944079216
        );
        
        core_inst_140097944079272: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944079272,
            fifo_full => fifo_full_140097944079272,
            outputs => outputs_140097944079272,
            outputs_full => outputs_full_140097944079272
        );
        
        core_inst_140097944079328: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944079328,
            fifo_full => fifo_full_140097944079328,
            outputs => outputs_140097944079328,
            outputs_full => outputs_full_140097944079328
        );
        
        core_inst_140097944079384: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944079384,
            fifo_full => fifo_full_140097944079384,
            outputs => outputs_140097944079384,
            outputs_full => outputs_full_140097944079384
        );
        
        core_inst_140097944079440: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944079440,
            fifo_full => fifo_full_140097944079440,
            outputs => outputs_140097944079440,
            outputs_full => outputs_full_140097944079440
        );
        
        core_inst_140097944079496: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944079496,
            fifo_full => fifo_full_140097944079496,
            outputs => outputs_140097944079496,
            outputs_full => outputs_full_140097944079496
        );
        
        core_inst_140097944079552: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944079552,
            fifo_full => fifo_full_140097944079552,
            outputs => outputs_140097944079552,
            outputs_full => outputs_full_140097944079552
        );
        
        core_inst_140097944079608: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944079608,
            fifo_full => fifo_full_140097944079608,
            outputs => outputs_140097944079608,
            outputs_full => outputs_full_140097944079608
        );
        
        core_inst_140097944079664: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944079664,
            fifo_full => fifo_full_140097944079664,
            outputs => outputs_140097944079664,
            outputs_full => outputs_full_140097944079664
        );
        
        core_inst_140097944079720: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944079720,
            fifo_full => fifo_full_140097944079720,
            outputs => outputs_140097944079720,
            outputs_full => outputs_full_140097944079720
        );
        
        core_inst_140097944079776: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944079776,
            fifo_full => fifo_full_140097944079776,
            outputs => outputs_140097944079776,
            outputs_full => outputs_full_140097944079776
        );
        
        core_inst_140097944079832: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944079832,
            fifo_full => fifo_full_140097944079832,
            outputs => outputs_140097944079832,
            outputs_full => outputs_full_140097944079832
        );
        
        core_inst_140097944079888: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944079888,
            fifo_full => fifo_full_140097944079888,
            outputs => outputs_140097944079888,
            outputs_full => outputs_full_140097944079888
        );
        
        core_inst_140097944079944: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944079944,
            fifo_full => fifo_full_140097944079944,
            outputs => outputs_140097944079944,
            outputs_full => outputs_full_140097944079944
        );
        
        core_inst_140097944080000: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944080000,
            fifo_full => fifo_full_140097944080000,
            outputs => outputs_140097944080000,
            outputs_full => outputs_full_140097944080000
        );
        
        core_inst_140097944080056: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944080056,
            fifo_full => fifo_full_140097944080056,
            outputs => outputs_140097944080056,
            outputs_full => outputs_full_140097944080056
        );
        
        core_inst_140097944080112: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944080112,
            fifo_full => fifo_full_140097944080112,
            outputs => outputs_140097944080112,
            outputs_full => outputs_full_140097944080112
        );
        
        core_inst_140097944080168: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944080168,
            fifo_full => fifo_full_140097944080168,
            outputs => outputs_140097944080168,
            outputs_full => outputs_full_140097944080168
        );
        
        core_inst_140097944080224: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944080224,
            fifo_full => fifo_full_140097944080224,
            outputs => outputs_140097944080224,
            outputs_full => outputs_full_140097944080224
        );
        
        core_inst_140097944080280: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944080280,
            fifo_full => fifo_full_140097944080280,
            outputs => outputs_140097944080280,
            outputs_full => outputs_full_140097944080280
        );
        
        core_inst_140097944080336: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944080336,
            fifo_full => fifo_full_140097944080336,
            outputs => outputs_140097944080336,
            outputs_full => outputs_full_140097944080336
        );
        
        core_inst_140097944096840: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944096840,
            fifo_full => fifo_full_140097944096840,
            outputs => outputs_140097944096840,
            outputs_full => outputs_full_140097944096840
        );
        
        core_inst_140097944096896: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944096896,
            fifo_full => fifo_full_140097944096896,
            outputs => outputs_140097944096896,
            outputs_full => outputs_full_140097944096896
        );
        
        core_inst_140097944096952: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944096952,
            fifo_full => fifo_full_140097944096952,
            outputs => outputs_140097944096952,
            outputs_full => outputs_full_140097944096952
        );
        
        core_inst_140097944097008: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944097008,
            fifo_full => fifo_full_140097944097008,
            outputs => outputs_140097944097008,
            outputs_full => outputs_full_140097944097008
        );
        
        core_inst_140097944097064: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944097064,
            fifo_full => fifo_full_140097944097064,
            outputs => outputs_140097944097064,
            outputs_full => outputs_full_140097944097064
        );
        
        core_inst_140097944097120: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944097120,
            fifo_full => fifo_full_140097944097120,
            outputs => outputs_140097944097120,
            outputs_full => outputs_full_140097944097120
        );
        
        core_inst_140097944097176: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944097176,
            fifo_full => fifo_full_140097944097176,
            outputs => outputs_140097944097176,
            outputs_full => outputs_full_140097944097176
        );
        
        core_inst_140097944097232: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944097232,
            fifo_full => fifo_full_140097944097232,
            outputs => outputs_140097944097232,
            outputs_full => outputs_full_140097944097232
        );
        
        core_inst_140097944097288: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944097288,
            fifo_full => fifo_full_140097944097288,
            outputs => outputs_140097944097288,
            outputs_full => outputs_full_140097944097288
        );
        
        core_inst_140097944097344: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944097344,
            fifo_full => fifo_full_140097944097344,
            outputs => outputs_140097944097344,
            outputs_full => outputs_full_140097944097344
        );
        
        core_inst_140097944097400: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944097400,
            fifo_full => fifo_full_140097944097400,
            outputs => outputs_140097944097400,
            outputs_full => outputs_full_140097944097400
        );
        
        core_inst_140097944097456: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944097456,
            fifo_full => fifo_full_140097944097456,
            outputs => outputs_140097944097456,
            outputs_full => outputs_full_140097944097456
        );
        
        core_inst_140097944097512: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944097512,
            fifo_full => fifo_full_140097944097512,
            outputs => outputs_140097944097512,
            outputs_full => outputs_full_140097944097512
        );
        
        core_inst_140097944097568: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944097568,
            fifo_full => fifo_full_140097944097568,
            outputs => outputs_140097944097568,
            outputs_full => outputs_full_140097944097568
        );
        
        core_inst_140097944097624: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944097624,
            fifo_full => fifo_full_140097944097624,
            outputs => outputs_140097944097624,
            outputs_full => outputs_full_140097944097624
        );
        
        core_inst_140097944097680: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944097680,
            fifo_full => fifo_full_140097944097680,
            outputs => outputs_140097944097680,
            outputs_full => outputs_full_140097944097680
        );
        
        core_inst_140097944097736: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944097736,
            fifo_full => fifo_full_140097944097736,
            outputs => outputs_140097944097736,
            outputs_full => outputs_full_140097944097736
        );
        
        core_inst_140097944097792: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944097792,
            fifo_full => fifo_full_140097944097792,
            outputs => outputs_140097944097792,
            outputs_full => outputs_full_140097944097792
        );
        
        core_inst_140097944097848: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944097848,
            fifo_full => fifo_full_140097944097848,
            outputs => outputs_140097944097848,
            outputs_full => outputs_full_140097944097848
        );
        
        core_inst_140097944097904: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944097904,
            fifo_full => fifo_full_140097944097904,
            outputs => outputs_140097944097904,
            outputs_full => outputs_full_140097944097904
        );
        
        core_inst_140097944097960: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944097960,
            fifo_full => fifo_full_140097944097960,
            outputs => outputs_140097944097960,
            outputs_full => outputs_full_140097944097960
        );
        
        core_inst_140097944098016: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944098016,
            fifo_full => fifo_full_140097944098016,
            outputs => outputs_140097944098016,
            outputs_full => outputs_full_140097944098016
        );
        
        core_inst_140097944098072: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944098072,
            fifo_full => fifo_full_140097944098072,
            outputs => outputs_140097944098072,
            outputs_full => outputs_full_140097944098072
        );
        
        core_inst_140097944098128: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944098128,
            fifo_full => fifo_full_140097944098128,
            outputs => outputs_140097944098128,
            outputs_full => outputs_full_140097944098128
        );
        
        core_inst_140097944098184: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944098184,
            fifo_full => fifo_full_140097944098184,
            outputs => outputs_140097944098184,
            outputs_full => outputs_full_140097944098184
        );
        
        core_inst_140097944098240: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944098240,
            fifo_full => fifo_full_140097944098240,
            outputs => outputs_140097944098240,
            outputs_full => outputs_full_140097944098240
        );
        
        core_inst_140097944098296: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944098296,
            fifo_full => fifo_full_140097944098296,
            outputs => outputs_140097944098296,
            outputs_full => outputs_full_140097944098296
        );
        
        core_inst_140097944098352: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944098352,
            fifo_full => fifo_full_140097944098352,
            outputs => outputs_140097944098352,
            outputs_full => outputs_full_140097944098352
        );
        
        core_inst_140097944098408: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944098408,
            fifo_full => fifo_full_140097944098408,
            outputs => outputs_140097944098408,
            outputs_full => outputs_full_140097944098408
        );
        
        core_inst_140097944098464: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944098464,
            fifo_full => fifo_full_140097944098464,
            outputs => outputs_140097944098464,
            outputs_full => outputs_full_140097944098464
        );
        
        core_inst_140097944098520: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944098520,
            fifo_full => fifo_full_140097944098520,
            outputs => outputs_140097944098520,
            outputs_full => outputs_full_140097944098520
        );
        
        core_inst_140097944098576: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944098576,
            fifo_full => fifo_full_140097944098576,
            outputs => outputs_140097944098576,
            outputs_full => outputs_full_140097944098576
        );
        
        core_inst_140097944098632: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944098632,
            fifo_full => fifo_full_140097944098632,
            outputs => outputs_140097944098632,
            outputs_full => outputs_full_140097944098632
        );
        
        core_inst_140097944098688: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944098688,
            fifo_full => fifo_full_140097944098688,
            outputs => outputs_140097944098688,
            outputs_full => outputs_full_140097944098688
        );
        
        core_inst_140097944098744: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944098744,
            fifo_full => fifo_full_140097944098744,
            outputs => outputs_140097944098744,
            outputs_full => outputs_full_140097944098744
        );
        
        core_inst_140097944098800: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944098800,
            fifo_full => fifo_full_140097944098800,
            outputs => outputs_140097944098800,
            outputs_full => outputs_full_140097944098800
        );
        
        core_inst_140097944098856: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944098856,
            fifo_full => fifo_full_140097944098856,
            outputs => outputs_140097944098856,
            outputs_full => outputs_full_140097944098856
        );
        
        core_inst_140097944098912: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944098912,
            fifo_full => fifo_full_140097944098912,
            outputs => outputs_140097944098912,
            outputs_full => outputs_full_140097944098912
        );
        
        core_inst_140097944098968: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944098968,
            fifo_full => fifo_full_140097944098968,
            outputs => outputs_140097944098968,
            outputs_full => outputs_full_140097944098968
        );
        
        core_inst_140097944099024: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944099024,
            fifo_full => fifo_full_140097944099024,
            outputs => outputs_140097944099024,
            outputs_full => outputs_full_140097944099024
        );
        
        core_inst_140097944099080: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944099080,
            fifo_full => fifo_full_140097944099080,
            outputs => outputs_140097944099080,
            outputs_full => outputs_full_140097944099080
        );
        
        core_inst_140097944099136: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944099136,
            fifo_full => fifo_full_140097944099136,
            outputs => outputs_140097944099136,
            outputs_full => outputs_full_140097944099136
        );
        
        core_inst_140097944099192: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944099192,
            fifo_full => fifo_full_140097944099192,
            outputs => outputs_140097944099192,
            outputs_full => outputs_full_140097944099192
        );
        
        core_inst_140097944099248: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944099248,
            fifo_full => fifo_full_140097944099248,
            outputs => outputs_140097944099248,
            outputs_full => outputs_full_140097944099248
        );
        
        core_inst_140097944099304: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944099304,
            fifo_full => fifo_full_140097944099304,
            outputs => outputs_140097944099304,
            outputs_full => outputs_full_140097944099304
        );
        
        core_inst_140097944099360: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944099360,
            fifo_full => fifo_full_140097944099360,
            outputs => outputs_140097944099360,
            outputs_full => outputs_full_140097944099360
        );
        
        core_inst_140097944099416: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944099416,
            fifo_full => fifo_full_140097944099416,
            outputs => outputs_140097944099416,
            outputs_full => outputs_full_140097944099416
        );
        
        core_inst_140097944099472: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944099472,
            fifo_full => fifo_full_140097944099472,
            outputs => outputs_140097944099472,
            outputs_full => outputs_full_140097944099472
        );
        
        core_inst_140097944099528: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944099528,
            fifo_full => fifo_full_140097944099528,
            outputs => outputs_140097944099528,
            outputs_full => outputs_full_140097944099528
        );
        
        core_inst_140097965543496: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097965543496,
            fifo_full => fifo_full_140097965543496,
            outputs => outputs_140097965543496,
            outputs_full => outputs_full_140097965543496
        );
        
        core_inst_140097944041736: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944041736,
            fifo_full => fifo_full_140097944041736,
            outputs => outputs_140097944041736,
            outputs_full => outputs_full_140097944041736
        );
        
        core_inst_140097944041624: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944041624,
            fifo_full => fifo_full_140097944041624,
            outputs => outputs_140097944041624,
            outputs_full => outputs_full_140097944041624
        );
        
        core_inst_140097944041568: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944041568,
            fifo_full => fifo_full_140097944041568,
            outputs => outputs_140097944041568,
            outputs_full => outputs_full_140097944041568
        );
        
        core_inst_140097944041792: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944041792,
            fifo_full => fifo_full_140097944041792,
            outputs => outputs_140097944041792,
            outputs_full => outputs_full_140097944041792
        );
        
        core_inst_140097944041456: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944041456,
            fifo_full => fifo_full_140097944041456,
            outputs => outputs_140097944041456,
            outputs_full => outputs_full_140097944041456
        );
        
        core_inst_140097944099584: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944099584,
            fifo_full => fifo_full_140097944099584,
            outputs => outputs_140097944099584,
            outputs_full => outputs_full_140097944099584
        );
        
        core_inst_140097944099640: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944099640,
            fifo_full => fifo_full_140097944099640,
            outputs => outputs_140097944099640,
            outputs_full => outputs_full_140097944099640
        );
        
        core_inst_140097944099696: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944099696,
            fifo_full => fifo_full_140097944099696,
            outputs => outputs_140097944099696,
            outputs_full => outputs_full_140097944099696
        );
        
        core_inst_140097944099752: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944099752,
            fifo_full => fifo_full_140097944099752,
            outputs => outputs_140097944099752,
            outputs_full => outputs_full_140097944099752
        );
        
        core_inst_140097944099808: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944099808,
            fifo_full => fifo_full_140097944099808,
            outputs => outputs_140097944099808,
            outputs_full => outputs_full_140097944099808
        );
        
        core_inst_140097944099864: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944099864,
            fifo_full => fifo_full_140097944099864,
            outputs => outputs_140097944099864,
            outputs_full => outputs_full_140097944099864
        );
        
        core_inst_140097944099920: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944099920,
            fifo_full => fifo_full_140097944099920,
            outputs => outputs_140097944099920,
            outputs_full => outputs_full_140097944099920
        );
        
        core_inst_140097944099976: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944099976,
            fifo_full => fifo_full_140097944099976,
            outputs => outputs_140097944099976,
            outputs_full => outputs_full_140097944099976
        );
        
        core_inst_140097944100032: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944100032,
            fifo_full => fifo_full_140097944100032,
            outputs => outputs_140097944100032,
            outputs_full => outputs_full_140097944100032
        );
        
        core_inst_140097944100088: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944100088,
            fifo_full => fifo_full_140097944100088,
            outputs => outputs_140097944100088,
            outputs_full => outputs_full_140097944100088
        );
        
        core_inst_140097944100144: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944100144,
            fifo_full => fifo_full_140097944100144,
            outputs => outputs_140097944100144,
            outputs_full => outputs_full_140097944100144
        );
        
        core_inst_140097944100200: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944100200,
            fifo_full => fifo_full_140097944100200,
            outputs => outputs_140097944100200,
            outputs_full => outputs_full_140097944100200
        );
        
        core_inst_140097944100256: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944100256,
            fifo_full => fifo_full_140097944100256,
            outputs => outputs_140097944100256,
            outputs_full => outputs_full_140097944100256
        );
        
        core_inst_140097944100312: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944100312,
            fifo_full => fifo_full_140097944100312,
            outputs => outputs_140097944100312,
            outputs_full => outputs_full_140097944100312
        );
        
        core_inst_140097944100368: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944100368,
            fifo_full => fifo_full_140097944100368,
            outputs => outputs_140097944100368,
            outputs_full => outputs_full_140097944100368
        );
        
        core_inst_140097944100424: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944100424,
            fifo_full => fifo_full_140097944100424,
            outputs => outputs_140097944100424,
            outputs_full => outputs_full_140097944100424
        );
        
        core_inst_140097944100480: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944100480,
            fifo_full => fifo_full_140097944100480,
            outputs => outputs_140097944100480,
            outputs_full => outputs_full_140097944100480
        );
        
        core_inst_140097944100536: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944100536,
            fifo_full => fifo_full_140097944100536,
            outputs => outputs_140097944100536,
            outputs_full => outputs_full_140097944100536
        );
        
        core_inst_140097944100592: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944100592,
            fifo_full => fifo_full_140097944100592,
            outputs => outputs_140097944100592,
            outputs_full => outputs_full_140097944100592
        );
        
        core_inst_140097944100648: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944100648,
            fifo_full => fifo_full_140097944100648,
            outputs => outputs_140097944100648,
            outputs_full => outputs_full_140097944100648
        );
        
        core_inst_140097944100704: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944100704,
            fifo_full => fifo_full_140097944100704,
            outputs => outputs_140097944100704,
            outputs_full => outputs_full_140097944100704
        );
        
        core_inst_140097944100760: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944100760,
            fifo_full => fifo_full_140097944100760,
            outputs => outputs_140097944100760,
            outputs_full => outputs_full_140097944100760
        );
        
        core_inst_140097944100816: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944100816,
            fifo_full => fifo_full_140097944100816,
            outputs => outputs_140097944100816,
            outputs_full => outputs_full_140097944100816
        );
        
        core_inst_140097944113224: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944113224,
            fifo_full => fifo_full_140097944113224,
            outputs => outputs_140097944113224,
            outputs_full => outputs_full_140097944113224
        );
        
        core_inst_140097944113280: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944113280,
            fifo_full => fifo_full_140097944113280,
            outputs => outputs_140097944113280,
            outputs_full => outputs_full_140097944113280
        );
        
        core_inst_140097944113336: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944113336,
            fifo_full => fifo_full_140097944113336,
            outputs => outputs_140097944113336,
            outputs_full => outputs_full_140097944113336
        );
        
        core_inst_140097944113392: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944113392,
            fifo_full => fifo_full_140097944113392,
            outputs => outputs_140097944113392,
            outputs_full => outputs_full_140097944113392
        );
        
        core_inst_140097944113448: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944113448,
            fifo_full => fifo_full_140097944113448,
            outputs => outputs_140097944113448,
            outputs_full => outputs_full_140097944113448
        );
        
        core_inst_140097944113504: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944113504,
            fifo_full => fifo_full_140097944113504,
            outputs => outputs_140097944113504,
            outputs_full => outputs_full_140097944113504
        );
        
        core_inst_140097944113560: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944113560,
            fifo_full => fifo_full_140097944113560,
            outputs => outputs_140097944113560,
            outputs_full => outputs_full_140097944113560
        );
        
        core_inst_140097944113616: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944113616,
            fifo_full => fifo_full_140097944113616,
            outputs => outputs_140097944113616,
            outputs_full => outputs_full_140097944113616
        );
        
        core_inst_140097944113672: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944113672,
            fifo_full => fifo_full_140097944113672,
            outputs => outputs_140097944113672,
            outputs_full => outputs_full_140097944113672
        );
        
        core_inst_140097944113728: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944113728,
            fifo_full => fifo_full_140097944113728,
            outputs => outputs_140097944113728,
            outputs_full => outputs_full_140097944113728
        );
        
        core_inst_140097944113784: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944113784,
            fifo_full => fifo_full_140097944113784,
            outputs => outputs_140097944113784,
            outputs_full => outputs_full_140097944113784
        );
        
        core_inst_140097944113840: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944113840,
            fifo_full => fifo_full_140097944113840,
            outputs => outputs_140097944113840,
            outputs_full => outputs_full_140097944113840
        );
        
        core_inst_140097944113896: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944113896,
            fifo_full => fifo_full_140097944113896,
            outputs => outputs_140097944113896,
            outputs_full => outputs_full_140097944113896
        );
        
        core_inst_140097944113952: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944113952,
            fifo_full => fifo_full_140097944113952,
            outputs => outputs_140097944113952,
            outputs_full => outputs_full_140097944113952
        );
        
        core_inst_140097944114008: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944114008,
            fifo_full => fifo_full_140097944114008,
            outputs => outputs_140097944114008,
            outputs_full => outputs_full_140097944114008
        );
        
        core_inst_140097944114064: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944114064,
            fifo_full => fifo_full_140097944114064,
            outputs => outputs_140097944114064,
            outputs_full => outputs_full_140097944114064
        );
        
        core_inst_140097944114120: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944114120,
            fifo_full => fifo_full_140097944114120,
            outputs => outputs_140097944114120,
            outputs_full => outputs_full_140097944114120
        );
        
        core_inst_140097944114176: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944114176,
            fifo_full => fifo_full_140097944114176,
            outputs => outputs_140097944114176,
            outputs_full => outputs_full_140097944114176
        );
        
        core_inst_140097944114232: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944114232,
            fifo_full => fifo_full_140097944114232,
            outputs => outputs_140097944114232,
            outputs_full => outputs_full_140097944114232
        );
        
        core_inst_140097944114288: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944114288,
            fifo_full => fifo_full_140097944114288,
            outputs => outputs_140097944114288,
            outputs_full => outputs_full_140097944114288
        );
        
        core_inst_140097944114344: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944114344,
            fifo_full => fifo_full_140097944114344,
            outputs => outputs_140097944114344,
            outputs_full => outputs_full_140097944114344
        );
        
        core_inst_140097944114400: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944114400,
            fifo_full => fifo_full_140097944114400,
            outputs => outputs_140097944114400,
            outputs_full => outputs_full_140097944114400
        );
        
        core_inst_140097944114456: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944114456,
            fifo_full => fifo_full_140097944114456,
            outputs => outputs_140097944114456,
            outputs_full => outputs_full_140097944114456
        );
        
        core_inst_140097944114512: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944114512,
            fifo_full => fifo_full_140097944114512,
            outputs => outputs_140097944114512,
            outputs_full => outputs_full_140097944114512
        );
        
        core_inst_140097944114568: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944114568,
            fifo_full => fifo_full_140097944114568,
            outputs => outputs_140097944114568,
            outputs_full => outputs_full_140097944114568
        );
        
        core_inst_140097944114624: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944114624,
            fifo_full => fifo_full_140097944114624,
            outputs => outputs_140097944114624,
            outputs_full => outputs_full_140097944114624
        );
        
        core_inst_140097944114680: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944114680,
            fifo_full => fifo_full_140097944114680,
            outputs => outputs_140097944114680,
            outputs_full => outputs_full_140097944114680
        );
        
        core_inst_140097944114736: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944114736,
            fifo_full => fifo_full_140097944114736,
            outputs => outputs_140097944114736,
            outputs_full => outputs_full_140097944114736
        );
        
        core_inst_140097944114792: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944114792,
            fifo_full => fifo_full_140097944114792,
            outputs => outputs_140097944114792,
            outputs_full => outputs_full_140097944114792
        );
        
        core_inst_140097944114848: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944114848,
            fifo_full => fifo_full_140097944114848,
            outputs => outputs_140097944114848,
            outputs_full => outputs_full_140097944114848
        );
        
        core_inst_140097944114904: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944114904,
            fifo_full => fifo_full_140097944114904,
            outputs => outputs_140097944114904,
            outputs_full => outputs_full_140097944114904
        );
        
        core_inst_140097944114960: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944114960,
            fifo_full => fifo_full_140097944114960,
            outputs => outputs_140097944114960,
            outputs_full => outputs_full_140097944114960
        );
        
        core_inst_140097944115016: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944115016,
            fifo_full => fifo_full_140097944115016,
            outputs => outputs_140097944115016,
            outputs_full => outputs_full_140097944115016
        );
        
        core_inst_140097944115072: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944115072,
            fifo_full => fifo_full_140097944115072,
            outputs => outputs_140097944115072,
            outputs_full => outputs_full_140097944115072
        );
        
        core_inst_140097944115128: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944115128,
            fifo_full => fifo_full_140097944115128,
            outputs => outputs_140097944115128,
            outputs_full => outputs_full_140097944115128
        );
        
        core_inst_140097944115184: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944115184,
            fifo_full => fifo_full_140097944115184,
            outputs => outputs_140097944115184,
            outputs_full => outputs_full_140097944115184
        );
        
        core_inst_140097944115240: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944115240,
            fifo_full => fifo_full_140097944115240,
            outputs => outputs_140097944115240,
            outputs_full => outputs_full_140097944115240
        );
        
        core_inst_140097944115296: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944115296,
            fifo_full => fifo_full_140097944115296,
            outputs => outputs_140097944115296,
            outputs_full => outputs_full_140097944115296
        );
        
        core_inst_140097944115352: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944115352,
            fifo_full => fifo_full_140097944115352,
            outputs => outputs_140097944115352,
            outputs_full => outputs_full_140097944115352
        );
        
        core_inst_140097944115408: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944115408,
            fifo_full => fifo_full_140097944115408,
            outputs => outputs_140097944115408,
            outputs_full => outputs_full_140097944115408
        );
        
        core_inst_140097944115464: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944115464,
            fifo_full => fifo_full_140097944115464,
            outputs => outputs_140097944115464,
            outputs_full => outputs_full_140097944115464
        );
        
        core_inst_140097944115520: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944115520,
            fifo_full => fifo_full_140097944115520,
            outputs => outputs_140097944115520,
            outputs_full => outputs_full_140097944115520
        );
        
        core_inst_140097944115576: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944115576,
            fifo_full => fifo_full_140097944115576,
            outputs => outputs_140097944115576,
            outputs_full => outputs_full_140097944115576
        );
        
        core_inst_140097944115632: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944115632,
            fifo_full => fifo_full_140097944115632,
            outputs => outputs_140097944115632,
            outputs_full => outputs_full_140097944115632
        );
        
        core_inst_140097944115688: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944115688,
            fifo_full => fifo_full_140097944115688,
            outputs => outputs_140097944115688,
            outputs_full => outputs_full_140097944115688
        );
        
        core_inst_140097944115744: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944115744,
            fifo_full => fifo_full_140097944115744,
            outputs => outputs_140097944115744,
            outputs_full => outputs_full_140097944115744
        );
        
        core_inst_140097944115800: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944115800,
            fifo_full => fifo_full_140097944115800,
            outputs => outputs_140097944115800,
            outputs_full => outputs_full_140097944115800
        );
        
        core_inst_140097944115856: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944115856,
            fifo_full => fifo_full_140097944115856,
            outputs => outputs_140097944115856,
            outputs_full => outputs_full_140097944115856
        );
        
        core_inst_140097944115912: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944115912,
            fifo_full => fifo_full_140097944115912,
            outputs => outputs_140097944115912,
            outputs_full => outputs_full_140097944115912
        );
        
        core_inst_140097944115968: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944115968,
            fifo_full => fifo_full_140097944115968,
            outputs => outputs_140097944115968,
            outputs_full => outputs_full_140097944115968
        );
        
        core_inst_140097944116024: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944116024,
            fifo_full => fifo_full_140097944116024,
            outputs => outputs_140097944116024,
            outputs_full => outputs_full_140097944116024
        );
        
        core_inst_140097944116080: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944116080,
            fifo_full => fifo_full_140097944116080,
            outputs => outputs_140097944116080,
            outputs_full => outputs_full_140097944116080
        );
        
        core_inst_140097944116136: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944116136,
            fifo_full => fifo_full_140097944116136,
            outputs => outputs_140097944116136,
            outputs_full => outputs_full_140097944116136
        );
        
        core_inst_140097944116192: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944116192,
            fifo_full => fifo_full_140097944116192,
            outputs => outputs_140097944116192,
            outputs_full => outputs_full_140097944116192
        );
        
        core_inst_140097944116248: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944116248,
            fifo_full => fifo_full_140097944116248,
            outputs => outputs_140097944116248,
            outputs_full => outputs_full_140097944116248
        );
        
        core_inst_140097944116304: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944116304,
            fifo_full => fifo_full_140097944116304,
            outputs => outputs_140097944116304,
            outputs_full => outputs_full_140097944116304
        );
        
        core_inst_140097944116360: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944116360,
            fifo_full => fifo_full_140097944116360,
            outputs => outputs_140097944116360,
            outputs_full => outputs_full_140097944116360
        );
        
        core_inst_140097944116416: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944116416,
            fifo_full => fifo_full_140097944116416,
            outputs => outputs_140097944116416,
            outputs_full => outputs_full_140097944116416
        );
        
        core_inst_140097944116472: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944116472,
            fifo_full => fifo_full_140097944116472,
            outputs => outputs_140097944116472,
            outputs_full => outputs_full_140097944116472
        );
        
        core_inst_140097944116528: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944116528,
            fifo_full => fifo_full_140097944116528,
            outputs => outputs_140097944116528,
            outputs_full => outputs_full_140097944116528
        );
        
        core_inst_140097944116584: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944116584,
            fifo_full => fifo_full_140097944116584,
            outputs => outputs_140097944116584,
            outputs_full => outputs_full_140097944116584
        );
        
        core_inst_140097944116640: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944116640,
            fifo_full => fifo_full_140097944116640,
            outputs => outputs_140097944116640,
            outputs_full => outputs_full_140097944116640
        );
        
        core_inst_140097944116696: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944116696,
            fifo_full => fifo_full_140097944116696,
            outputs => outputs_140097944116696,
            outputs_full => outputs_full_140097944116696
        );
        
        core_inst_140097944116752: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944116752,
            fifo_full => fifo_full_140097944116752,
            outputs => outputs_140097944116752,
            outputs_full => outputs_full_140097944116752
        );
        
        core_inst_140097944116808: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944116808,
            fifo_full => fifo_full_140097944116808,
            outputs => outputs_140097944116808,
            outputs_full => outputs_full_140097944116808
        );
        
        core_inst_140097944116864: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944116864,
            fifo_full => fifo_full_140097944116864,
            outputs => outputs_140097944116864,
            outputs_full => outputs_full_140097944116864
        );
        
        core_inst_140097944116920: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944116920,
            fifo_full => fifo_full_140097944116920,
            outputs => outputs_140097944116920,
            outputs_full => outputs_full_140097944116920
        );
        
        core_inst_140097944116976: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944116976,
            fifo_full => fifo_full_140097944116976,
            outputs => outputs_140097944116976,
            outputs_full => outputs_full_140097944116976
        );
        
        core_inst_140097944117032: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944117032,
            fifo_full => fifo_full_140097944117032,
            outputs => outputs_140097944117032,
            outputs_full => outputs_full_140097944117032
        );
        
        core_inst_140097944117088: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944117088,
            fifo_full => fifo_full_140097944117088,
            outputs => outputs_140097944117088,
            outputs_full => outputs_full_140097944117088
        );
        
        core_inst_140097944117144: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944117144,
            fifo_full => fifo_full_140097944117144,
            outputs => outputs_140097944117144,
            outputs_full => outputs_full_140097944117144
        );
        
        core_inst_140097944117200: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944117200,
            fifo_full => fifo_full_140097944117200,
            outputs => outputs_140097944117200,
            outputs_full => outputs_full_140097944117200
        );
        
        core_inst_140097944125512: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944125512,
            fifo_full => fifo_full_140097944125512,
            outputs => outputs_140097944125512,
            outputs_full => outputs_full_140097944125512
        );
        
        core_inst_140097944125568: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944125568,
            fifo_full => fifo_full_140097944125568,
            outputs => outputs_140097944125568,
            outputs_full => outputs_full_140097944125568
        );
        
        core_inst_140097944125624: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944125624,
            fifo_full => fifo_full_140097944125624,
            outputs => outputs_140097944125624,
            outputs_full => outputs_full_140097944125624
        );
        
        core_inst_140097944125680: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944125680,
            fifo_full => fifo_full_140097944125680,
            outputs => outputs_140097944125680,
            outputs_full => outputs_full_140097944125680
        );
        
        core_inst_140097944125736: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944125736,
            fifo_full => fifo_full_140097944125736,
            outputs => outputs_140097944125736,
            outputs_full => outputs_full_140097944125736
        );
        
        core_inst_140097944125792: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944125792,
            fifo_full => fifo_full_140097944125792,
            outputs => outputs_140097944125792,
            outputs_full => outputs_full_140097944125792
        );
        
        core_inst_140097944125848: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944125848,
            fifo_full => fifo_full_140097944125848,
            outputs => outputs_140097944125848,
            outputs_full => outputs_full_140097944125848
        );
        
        core_inst_140097944125904: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944125904,
            fifo_full => fifo_full_140097944125904,
            outputs => outputs_140097944125904,
            outputs_full => outputs_full_140097944125904
        );
        
        core_inst_140097944125960: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944125960,
            fifo_full => fifo_full_140097944125960,
            outputs => outputs_140097944125960,
            outputs_full => outputs_full_140097944125960
        );
        
        core_inst_140097944126016: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944126016,
            fifo_full => fifo_full_140097944126016,
            outputs => outputs_140097944126016,
            outputs_full => outputs_full_140097944126016
        );
        
        core_inst_140097944126072: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944126072,
            fifo_full => fifo_full_140097944126072,
            outputs => outputs_140097944126072,
            outputs_full => outputs_full_140097944126072
        );
        
        core_inst_140097944126128: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944126128,
            fifo_full => fifo_full_140097944126128,
            outputs => outputs_140097944126128,
            outputs_full => outputs_full_140097944126128
        );
        
        core_inst_140097944126184: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944126184,
            fifo_full => fifo_full_140097944126184,
            outputs => outputs_140097944126184,
            outputs_full => outputs_full_140097944126184
        );
        
        core_inst_140097944126240: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944126240,
            fifo_full => fifo_full_140097944126240,
            outputs => outputs_140097944126240,
            outputs_full => outputs_full_140097944126240
        );
        
        core_inst_140097944126296: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944126296,
            fifo_full => fifo_full_140097944126296,
            outputs => outputs_140097944126296,
            outputs_full => outputs_full_140097944126296
        );
        
        core_inst_140097944126352: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944126352,
            fifo_full => fifo_full_140097944126352,
            outputs => outputs_140097944126352,
            outputs_full => outputs_full_140097944126352
        );
        
        core_inst_140097944126408: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944126408,
            fifo_full => fifo_full_140097944126408,
            outputs => outputs_140097944126408,
            outputs_full => outputs_full_140097944126408
        );
        
        core_inst_140097944126464: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944126464,
            fifo_full => fifo_full_140097944126464,
            outputs => outputs_140097944126464,
            outputs_full => outputs_full_140097944126464
        );
        
        core_inst_140097944126520: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944126520,
            fifo_full => fifo_full_140097944126520,
            outputs => outputs_140097944126520,
            outputs_full => outputs_full_140097944126520
        );
        
        core_inst_140097944126576: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944126576,
            fifo_full => fifo_full_140097944126576,
            outputs => outputs_140097944126576,
            outputs_full => outputs_full_140097944126576
        );
        
        core_inst_140097944126632: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944126632,
            fifo_full => fifo_full_140097944126632,
            outputs => outputs_140097944126632,
            outputs_full => outputs_full_140097944126632
        );
        
        core_inst_140097944126688: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944126688,
            fifo_full => fifo_full_140097944126688,
            outputs => outputs_140097944126688,
            outputs_full => outputs_full_140097944126688
        );
        
        core_inst_140097944126744: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944126744,
            fifo_full => fifo_full_140097944126744,
            outputs => outputs_140097944126744,
            outputs_full => outputs_full_140097944126744
        );
        
        core_inst_140097944126800: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944126800,
            fifo_full => fifo_full_140097944126800,
            outputs => outputs_140097944126800,
            outputs_full => outputs_full_140097944126800
        );
        
        core_inst_140097944126856: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944126856,
            fifo_full => fifo_full_140097944126856,
            outputs => outputs_140097944126856,
            outputs_full => outputs_full_140097944126856
        );
        
        core_inst_140097944126912: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944126912,
            fifo_full => fifo_full_140097944126912,
            outputs => outputs_140097944126912,
            outputs_full => outputs_full_140097944126912
        );
        
        core_inst_140097944126968: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944126968,
            fifo_full => fifo_full_140097944126968,
            outputs => outputs_140097944126968,
            outputs_full => outputs_full_140097944126968
        );
        
        core_inst_140097944127024: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944127024,
            fifo_full => fifo_full_140097944127024,
            outputs => outputs_140097944127024,
            outputs_full => outputs_full_140097944127024
        );
        
        core_inst_140097944127080: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944127080,
            fifo_full => fifo_full_140097944127080,
            outputs => outputs_140097944127080,
            outputs_full => outputs_full_140097944127080
        );
        
        core_inst_140097944127136: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944127136,
            fifo_full => fifo_full_140097944127136,
            outputs => outputs_140097944127136,
            outputs_full => outputs_full_140097944127136
        );
        
        core_inst_140097944127192: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944127192,
            fifo_full => fifo_full_140097944127192,
            outputs => outputs_140097944127192,
            outputs_full => outputs_full_140097944127192
        );
        
        core_inst_140097944127248: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944127248,
            fifo_full => fifo_full_140097944127248,
            outputs => outputs_140097944127248,
            outputs_full => outputs_full_140097944127248
        );
        
        core_inst_140097944127304: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944127304,
            fifo_full => fifo_full_140097944127304,
            outputs => outputs_140097944127304,
            outputs_full => outputs_full_140097944127304
        );
        
        core_inst_140097944127360: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944127360,
            fifo_full => fifo_full_140097944127360,
            outputs => outputs_140097944127360,
            outputs_full => outputs_full_140097944127360
        );
        
        core_inst_140097944127416: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944127416,
            fifo_full => fifo_full_140097944127416,
            outputs => outputs_140097944127416,
            outputs_full => outputs_full_140097944127416
        );
        
        core_inst_140097944127472: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944127472,
            fifo_full => fifo_full_140097944127472,
            outputs => outputs_140097944127472,
            outputs_full => outputs_full_140097944127472
        );
        
        core_inst_140097944127528: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944127528,
            fifo_full => fifo_full_140097944127528,
            outputs => outputs_140097944127528,
            outputs_full => outputs_full_140097944127528
        );
        
        core_inst_140097944127584: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944127584,
            fifo_full => fifo_full_140097944127584,
            outputs => outputs_140097944127584,
            outputs_full => outputs_full_140097944127584
        );
        
        core_inst_140097944127640: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944127640,
            fifo_full => fifo_full_140097944127640,
            outputs => outputs_140097944127640,
            outputs_full => outputs_full_140097944127640
        );
        
        core_inst_140097944127696: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944127696,
            fifo_full => fifo_full_140097944127696,
            outputs => outputs_140097944127696,
            outputs_full => outputs_full_140097944127696
        );
        
        core_inst_140097944127752: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944127752,
            fifo_full => fifo_full_140097944127752,
            outputs => outputs_140097944127752,
            outputs_full => outputs_full_140097944127752
        );
        
        core_inst_140097944127808: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944127808,
            fifo_full => fifo_full_140097944127808,
            outputs => outputs_140097944127808,
            outputs_full => outputs_full_140097944127808
        );
        
        core_inst_140097944127864: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944127864,
            fifo_full => fifo_full_140097944127864,
            outputs => outputs_140097944127864,
            outputs_full => outputs_full_140097944127864
        );
        
        core_inst_140097944127920: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944127920,
            fifo_full => fifo_full_140097944127920,
            outputs => outputs_140097944127920,
            outputs_full => outputs_full_140097944127920
        );
        
        core_inst_140097944127976: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944127976,
            fifo_full => fifo_full_140097944127976,
            outputs => outputs_140097944127976,
            outputs_full => outputs_full_140097944127976
        );
        
        core_inst_140097944128032: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944128032,
            fifo_full => fifo_full_140097944128032,
            outputs => outputs_140097944128032,
            outputs_full => outputs_full_140097944128032
        );
        
        core_inst_140097944128088: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944128088,
            fifo_full => fifo_full_140097944128088,
            outputs => outputs_140097944128088,
            outputs_full => outputs_full_140097944128088
        );
        
        core_inst_140097944128144: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944128144,
            fifo_full => fifo_full_140097944128144,
            outputs => outputs_140097944128144,
            outputs_full => outputs_full_140097944128144
        );
        
        core_inst_140097944128200: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944128200,
            fifo_full => fifo_full_140097944128200,
            outputs => outputs_140097944128200,
            outputs_full => outputs_full_140097944128200
        );
        
        core_inst_140097944128256: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944128256,
            fifo_full => fifo_full_140097944128256,
            outputs => outputs_140097944128256,
            outputs_full => outputs_full_140097944128256
        );
        
        core_inst_140097944128312: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944128312,
            fifo_full => fifo_full_140097944128312,
            outputs => outputs_140097944128312,
            outputs_full => outputs_full_140097944128312
        );
        
        core_inst_140097944128368: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944128368,
            fifo_full => fifo_full_140097944128368,
            outputs => outputs_140097944128368,
            outputs_full => outputs_full_140097944128368
        );
        
        core_inst_140097944128424: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944128424,
            fifo_full => fifo_full_140097944128424,
            outputs => outputs_140097944128424,
            outputs_full => outputs_full_140097944128424
        );
        
        core_inst_140097944128480: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944128480,
            fifo_full => fifo_full_140097944128480,
            outputs => outputs_140097944128480,
            outputs_full => outputs_full_140097944128480
        );
        
        core_inst_140097944128536: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944128536,
            fifo_full => fifo_full_140097944128536,
            outputs => outputs_140097944128536,
            outputs_full => outputs_full_140097944128536
        );
        
        core_inst_140097944128592: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944128592,
            fifo_full => fifo_full_140097944128592,
            outputs => outputs_140097944128592,
            outputs_full => outputs_full_140097944128592
        );
        
        core_inst_140097944128648: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944128648,
            fifo_full => fifo_full_140097944128648,
            outputs => outputs_140097944128648,
            outputs_full => outputs_full_140097944128648
        );
        
        core_inst_140097944128704: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944128704,
            fifo_full => fifo_full_140097944128704,
            outputs => outputs_140097944128704,
            outputs_full => outputs_full_140097944128704
        );
        
        core_inst_140097944128760: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944128760,
            fifo_full => fifo_full_140097944128760,
            outputs => outputs_140097944128760,
            outputs_full => outputs_full_140097944128760
        );
        
        core_inst_140097944128816: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944128816,
            fifo_full => fifo_full_140097944128816,
            outputs => outputs_140097944128816,
            outputs_full => outputs_full_140097944128816
        );
        
        core_inst_140097944128872: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944128872,
            fifo_full => fifo_full_140097944128872,
            outputs => outputs_140097944128872,
            outputs_full => outputs_full_140097944128872
        );
        
        core_inst_140097944128928: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944128928,
            fifo_full => fifo_full_140097944128928,
            outputs => outputs_140097944128928,
            outputs_full => outputs_full_140097944128928
        );
        
        core_inst_140097944128984: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944128984,
            fifo_full => fifo_full_140097944128984,
            outputs => outputs_140097944128984,
            outputs_full => outputs_full_140097944128984
        );
        
        core_inst_140097944129040: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944129040,
            fifo_full => fifo_full_140097944129040,
            outputs => outputs_140097944129040,
            outputs_full => outputs_full_140097944129040
        );
        
        core_inst_140097944129096: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944129096,
            fifo_full => fifo_full_140097944129096,
            outputs => outputs_140097944129096,
            outputs_full => outputs_full_140097944129096
        );
        
        core_inst_140097944129152: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944129152,
            fifo_full => fifo_full_140097944129152,
            outputs => outputs_140097944129152,
            outputs_full => outputs_full_140097944129152
        );
        
        core_inst_140097944129208: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944129208,
            fifo_full => fifo_full_140097944129208,
            outputs => outputs_140097944129208,
            outputs_full => outputs_full_140097944129208
        );
        
        core_inst_140097944129264: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944129264,
            fifo_full => fifo_full_140097944129264,
            outputs => outputs_140097944129264,
            outputs_full => outputs_full_140097944129264
        );
        
        core_inst_140097944129320: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944129320,
            fifo_full => fifo_full_140097944129320,
            outputs => outputs_140097944129320,
            outputs_full => outputs_full_140097944129320
        );
        
        core_inst_140097944129376: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944129376,
            fifo_full => fifo_full_140097944129376,
            outputs => outputs_140097944129376,
            outputs_full => outputs_full_140097944129376
        );
        
        core_inst_140097944129432: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944129432,
            fifo_full => fifo_full_140097944129432,
            outputs => outputs_140097944129432,
            outputs_full => outputs_full_140097944129432
        );
        
        core_inst_140097944129488: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944129488,
            fifo_full => fifo_full_140097944129488,
            outputs => outputs_140097944129488,
            outputs_full => outputs_full_140097944129488
        );
        
        core_inst_140097944141896: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944141896,
            fifo_full => fifo_full_140097944141896,
            outputs => outputs_140097944141896,
            outputs_full => outputs_full_140097944141896
        );
        
        core_inst_140097944141952: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944141952,
            fifo_full => fifo_full_140097944141952,
            outputs => outputs_140097944141952,
            outputs_full => outputs_full_140097944141952
        );
        
        core_inst_140097944142008: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944142008,
            fifo_full => fifo_full_140097944142008,
            outputs => outputs_140097944142008,
            outputs_full => outputs_full_140097944142008
        );
        
        core_inst_140097944142064: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944142064,
            fifo_full => fifo_full_140097944142064,
            outputs => outputs_140097944142064,
            outputs_full => outputs_full_140097944142064
        );
        
        core_inst_140097944142120: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944142120,
            fifo_full => fifo_full_140097944142120,
            outputs => outputs_140097944142120,
            outputs_full => outputs_full_140097944142120
        );
        
        core_inst_140097944142176: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944142176,
            fifo_full => fifo_full_140097944142176,
            outputs => outputs_140097944142176,
            outputs_full => outputs_full_140097944142176
        );
        
        core_inst_140097944142232: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944142232,
            fifo_full => fifo_full_140097944142232,
            outputs => outputs_140097944142232,
            outputs_full => outputs_full_140097944142232
        );
        
        core_inst_140097944142288: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944142288,
            fifo_full => fifo_full_140097944142288,
            outputs => outputs_140097944142288,
            outputs_full => outputs_full_140097944142288
        );
        
        core_inst_140097944142344: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944142344,
            fifo_full => fifo_full_140097944142344,
            outputs => outputs_140097944142344,
            outputs_full => outputs_full_140097944142344
        );
        
        core_inst_140097944142400: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944142400,
            fifo_full => fifo_full_140097944142400,
            outputs => outputs_140097944142400,
            outputs_full => outputs_full_140097944142400
        );
        
        core_inst_140097944142456: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944142456,
            fifo_full => fifo_full_140097944142456,
            outputs => outputs_140097944142456,
            outputs_full => outputs_full_140097944142456
        );
        
        core_inst_140097944142512: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944142512,
            fifo_full => fifo_full_140097944142512,
            outputs => outputs_140097944142512,
            outputs_full => outputs_full_140097944142512
        );
        
        core_inst_140097944142568: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944142568,
            fifo_full => fifo_full_140097944142568,
            outputs => outputs_140097944142568,
            outputs_full => outputs_full_140097944142568
        );
        
        core_inst_140097944142624: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944142624,
            fifo_full => fifo_full_140097944142624,
            outputs => outputs_140097944142624,
            outputs_full => outputs_full_140097944142624
        );
        
        core_inst_140097944142680: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944142680,
            fifo_full => fifo_full_140097944142680,
            outputs => outputs_140097944142680,
            outputs_full => outputs_full_140097944142680
        );
        
        core_inst_140097944142736: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944142736,
            fifo_full => fifo_full_140097944142736,
            outputs => outputs_140097944142736,
            outputs_full => outputs_full_140097944142736
        );
        
        core_inst_140097944142792: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944142792,
            fifo_full => fifo_full_140097944142792,
            outputs => outputs_140097944142792,
            outputs_full => outputs_full_140097944142792
        );
        
        core_inst_140097944142848: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944142848,
            fifo_full => fifo_full_140097944142848,
            outputs => outputs_140097944142848,
            outputs_full => outputs_full_140097944142848
        );
        
        core_inst_140097944142904: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944142904,
            fifo_full => fifo_full_140097944142904,
            outputs => outputs_140097944142904,
            outputs_full => outputs_full_140097944142904
        );
        
        core_inst_140097944142960: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944142960,
            fifo_full => fifo_full_140097944142960,
            outputs => outputs_140097944142960,
            outputs_full => outputs_full_140097944142960
        );
        
        core_inst_140097944143016: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944143016,
            fifo_full => fifo_full_140097944143016,
            outputs => outputs_140097944143016,
            outputs_full => outputs_full_140097944143016
        );
        
        core_inst_140097944143072: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944143072,
            fifo_full => fifo_full_140097944143072,
            outputs => outputs_140097944143072,
            outputs_full => outputs_full_140097944143072
        );
        
        core_inst_140097944143128: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944143128,
            fifo_full => fifo_full_140097944143128,
            outputs => outputs_140097944143128,
            outputs_full => outputs_full_140097944143128
        );
        
        core_inst_140097944143184: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944143184,
            fifo_full => fifo_full_140097944143184,
            outputs => outputs_140097944143184,
            outputs_full => outputs_full_140097944143184
        );
        
        core_inst_140097944143240: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944143240,
            fifo_full => fifo_full_140097944143240,
            outputs => outputs_140097944143240,
            outputs_full => outputs_full_140097944143240
        );
        
        core_inst_140097944143296: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944143296,
            fifo_full => fifo_full_140097944143296,
            outputs => outputs_140097944143296,
            outputs_full => outputs_full_140097944143296
        );
        
        core_inst_140097944143352: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944143352,
            fifo_full => fifo_full_140097944143352,
            outputs => outputs_140097944143352,
            outputs_full => outputs_full_140097944143352
        );
        
        core_inst_140097944143408: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944143408,
            fifo_full => fifo_full_140097944143408,
            outputs => outputs_140097944143408,
            outputs_full => outputs_full_140097944143408
        );
        
        core_inst_140097944143464: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944143464,
            fifo_full => fifo_full_140097944143464,
            outputs => outputs_140097944143464,
            outputs_full => outputs_full_140097944143464
        );
        
        core_inst_140097944143520: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944143520,
            fifo_full => fifo_full_140097944143520,
            outputs => outputs_140097944143520,
            outputs_full => outputs_full_140097944143520
        );
        
        core_inst_140097944143576: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944143576,
            fifo_full => fifo_full_140097944143576,
            outputs => outputs_140097944143576,
            outputs_full => outputs_full_140097944143576
        );
        
        core_inst_140097944143632: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944143632,
            fifo_full => fifo_full_140097944143632,
            outputs => outputs_140097944143632,
            outputs_full => outputs_full_140097944143632
        );
        
        core_inst_140097944143688: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944143688,
            fifo_full => fifo_full_140097944143688,
            outputs => outputs_140097944143688,
            outputs_full => outputs_full_140097944143688
        );
        
        core_inst_140097944143744: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944143744,
            fifo_full => fifo_full_140097944143744,
            outputs => outputs_140097944143744,
            outputs_full => outputs_full_140097944143744
        );
        
        core_inst_140097944143800: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944143800,
            fifo_full => fifo_full_140097944143800,
            outputs => outputs_140097944143800,
            outputs_full => outputs_full_140097944143800
        );
        
        core_inst_140097944143856: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944143856,
            fifo_full => fifo_full_140097944143856,
            outputs => outputs_140097944143856,
            outputs_full => outputs_full_140097944143856
        );
        
        core_inst_140097944143912: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944143912,
            fifo_full => fifo_full_140097944143912,
            outputs => outputs_140097944143912,
            outputs_full => outputs_full_140097944143912
        );
        
        core_inst_140097944143968: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944143968,
            fifo_full => fifo_full_140097944143968,
            outputs => outputs_140097944143968,
            outputs_full => outputs_full_140097944143968
        );
        
        core_inst_140097944144024: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944144024,
            fifo_full => fifo_full_140097944144024,
            outputs => outputs_140097944144024,
            outputs_full => outputs_full_140097944144024
        );
        
        core_inst_140097944144080: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944144080,
            fifo_full => fifo_full_140097944144080,
            outputs => outputs_140097944144080,
            outputs_full => outputs_full_140097944144080
        );
        
        core_inst_140097944144136: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944144136,
            fifo_full => fifo_full_140097944144136,
            outputs => outputs_140097944144136,
            outputs_full => outputs_full_140097944144136
        );
        
        core_inst_140097944144192: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944144192,
            fifo_full => fifo_full_140097944144192,
            outputs => outputs_140097944144192,
            outputs_full => outputs_full_140097944144192
        );
        
        core_inst_140097944144248: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944144248,
            fifo_full => fifo_full_140097944144248,
            outputs => outputs_140097944144248,
            outputs_full => outputs_full_140097944144248
        );
        
        core_inst_140097944144304: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944144304,
            fifo_full => fifo_full_140097944144304,
            outputs => outputs_140097944144304,
            outputs_full => outputs_full_140097944144304
        );
        
        core_inst_140097944144360: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944144360,
            fifo_full => fifo_full_140097944144360,
            outputs => outputs_140097944144360,
            outputs_full => outputs_full_140097944144360
        );
        
        core_inst_140097944144416: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944144416,
            fifo_full => fifo_full_140097944144416,
            outputs => outputs_140097944144416,
            outputs_full => outputs_full_140097944144416
        );
        
        core_inst_140097944144472: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944144472,
            fifo_full => fifo_full_140097944144472,
            outputs => outputs_140097944144472,
            outputs_full => outputs_full_140097944144472
        );
        
        core_inst_140097944144528: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944144528,
            fifo_full => fifo_full_140097944144528,
            outputs => outputs_140097944144528,
            outputs_full => outputs_full_140097944144528
        );
        
        core_inst_140097944144584: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944144584,
            fifo_full => fifo_full_140097944144584,
            outputs => outputs_140097944144584,
            outputs_full => outputs_full_140097944144584
        );
        
        core_inst_140097944144640: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944144640,
            fifo_full => fifo_full_140097944144640,
            outputs => outputs_140097944144640,
            outputs_full => outputs_full_140097944144640
        );
        
        core_inst_140097944144696: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944144696,
            fifo_full => fifo_full_140097944144696,
            outputs => outputs_140097944144696,
            outputs_full => outputs_full_140097944144696
        );
        
        core_inst_140097944144752: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944144752,
            fifo_full => fifo_full_140097944144752,
            outputs => outputs_140097944144752,
            outputs_full => outputs_full_140097944144752
        );
        
        core_inst_140097944144808: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944144808,
            fifo_full => fifo_full_140097944144808,
            outputs => outputs_140097944144808,
            outputs_full => outputs_full_140097944144808
        );
        
        core_inst_140097944144864: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944144864,
            fifo_full => fifo_full_140097944144864,
            outputs => outputs_140097944144864,
            outputs_full => outputs_full_140097944144864
        );
        
        core_inst_140097944144920: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944144920,
            fifo_full => fifo_full_140097944144920,
            outputs => outputs_140097944144920,
            outputs_full => outputs_full_140097944144920
        );
        
        core_inst_140097944144976: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944144976,
            fifo_full => fifo_full_140097944144976,
            outputs => outputs_140097944144976,
            outputs_full => outputs_full_140097944144976
        );
        
        core_inst_140097944145032: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944145032,
            fifo_full => fifo_full_140097944145032,
            outputs => outputs_140097944145032,
            outputs_full => outputs_full_140097944145032
        );
        
        core_inst_140097944145088: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944145088,
            fifo_full => fifo_full_140097944145088,
            outputs => outputs_140097944145088,
            outputs_full => outputs_full_140097944145088
        );
        
        core_inst_140097944145144: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944145144,
            fifo_full => fifo_full_140097944145144,
            outputs => outputs_140097944145144,
            outputs_full => outputs_full_140097944145144
        );
        
        core_inst_140097944145200: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944145200,
            fifo_full => fifo_full_140097944145200,
            outputs => outputs_140097944145200,
            outputs_full => outputs_full_140097944145200
        );
        
        core_inst_140097944145256: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944145256,
            fifo_full => fifo_full_140097944145256,
            outputs => outputs_140097944145256,
            outputs_full => outputs_full_140097944145256
        );
        
        core_inst_140097944145312: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944145312,
            fifo_full => fifo_full_140097944145312,
            outputs => outputs_140097944145312,
            outputs_full => outputs_full_140097944145312
        );
        
        core_inst_140097944145368: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944145368,
            fifo_full => fifo_full_140097944145368,
            outputs => outputs_140097944145368,
            outputs_full => outputs_full_140097944145368
        );
        
        core_inst_140097944145424: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944145424,
            fifo_full => fifo_full_140097944145424,
            outputs => outputs_140097944145424,
            outputs_full => outputs_full_140097944145424
        );
        
        core_inst_140097944145480: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944145480,
            fifo_full => fifo_full_140097944145480,
            outputs => outputs_140097944145480,
            outputs_full => outputs_full_140097944145480
        );
        
        core_inst_140097944145536: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944145536,
            fifo_full => fifo_full_140097944145536,
            outputs => outputs_140097944145536,
            outputs_full => outputs_full_140097944145536
        );
        
        core_inst_140097944145592: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944145592,
            fifo_full => fifo_full_140097944145592,
            outputs => outputs_140097944145592,
            outputs_full => outputs_full_140097944145592
        );
        
        core_inst_140097944145648: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944145648,
            fifo_full => fifo_full_140097944145648,
            outputs => outputs_140097944145648,
            outputs_full => outputs_full_140097944145648
        );
        
        core_inst_140097944145704: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944145704,
            fifo_full => fifo_full_140097944145704,
            outputs => outputs_140097944145704,
            outputs_full => outputs_full_140097944145704
        );
        
        core_inst_140097944145760: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944145760,
            fifo_full => fifo_full_140097944145760,
            outputs => outputs_140097944145760,
            outputs_full => outputs_full_140097944145760
        );
        
        core_inst_140097944145816: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944145816,
            fifo_full => fifo_full_140097944145816,
            outputs => outputs_140097944145816,
            outputs_full => outputs_full_140097944145816
        );
        
        core_inst_140097944145872: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944145872,
            fifo_full => fifo_full_140097944145872,
            outputs => outputs_140097944145872,
            outputs_full => outputs_full_140097944145872
        );
        
        core_inst_140097944154184: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944154184,
            fifo_full => fifo_full_140097944154184,
            outputs => outputs_140097944154184,
            outputs_full => outputs_full_140097944154184
        );
        
        core_inst_140097944154240: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944154240,
            fifo_full => fifo_full_140097944154240,
            outputs => outputs_140097944154240,
            outputs_full => outputs_full_140097944154240
        );
        
        core_inst_140097944154296: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944154296,
            fifo_full => fifo_full_140097944154296,
            outputs => outputs_140097944154296,
            outputs_full => outputs_full_140097944154296
        );
        
        core_inst_140097944154352: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944154352,
            fifo_full => fifo_full_140097944154352,
            outputs => outputs_140097944154352,
            outputs_full => outputs_full_140097944154352
        );
        
        core_inst_140097944154408: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944154408,
            fifo_full => fifo_full_140097944154408,
            outputs => outputs_140097944154408,
            outputs_full => outputs_full_140097944154408
        );
        
        core_inst_140097944154464: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944154464,
            fifo_full => fifo_full_140097944154464,
            outputs => outputs_140097944154464,
            outputs_full => outputs_full_140097944154464
        );
        
        core_inst_140097944154520: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944154520,
            fifo_full => fifo_full_140097944154520,
            outputs => outputs_140097944154520,
            outputs_full => outputs_full_140097944154520
        );
        
        core_inst_140097944154576: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944154576,
            fifo_full => fifo_full_140097944154576,
            outputs => outputs_140097944154576,
            outputs_full => outputs_full_140097944154576
        );
        
        core_inst_140097944154632: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944154632,
            fifo_full => fifo_full_140097944154632,
            outputs => outputs_140097944154632,
            outputs_full => outputs_full_140097944154632
        );
        
        core_inst_140097944154688: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944154688,
            fifo_full => fifo_full_140097944154688,
            outputs => outputs_140097944154688,
            outputs_full => outputs_full_140097944154688
        );
        
        core_inst_140097944154744: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944154744,
            fifo_full => fifo_full_140097944154744,
            outputs => outputs_140097944154744,
            outputs_full => outputs_full_140097944154744
        );
        
        core_inst_140097944154800: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944154800,
            fifo_full => fifo_full_140097944154800,
            outputs => outputs_140097944154800,
            outputs_full => outputs_full_140097944154800
        );
        
        core_inst_140097944154856: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944154856,
            fifo_full => fifo_full_140097944154856,
            outputs => outputs_140097944154856,
            outputs_full => outputs_full_140097944154856
        );
        
        core_inst_140097944154912: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944154912,
            fifo_full => fifo_full_140097944154912,
            outputs => outputs_140097944154912,
            outputs_full => outputs_full_140097944154912
        );
        
        core_inst_140097944154968: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944154968,
            fifo_full => fifo_full_140097944154968,
            outputs => outputs_140097944154968,
            outputs_full => outputs_full_140097944154968
        );
        
        core_inst_140097944155024: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944155024,
            fifo_full => fifo_full_140097944155024,
            outputs => outputs_140097944155024,
            outputs_full => outputs_full_140097944155024
        );
        
        core_inst_140097944155080: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944155080,
            fifo_full => fifo_full_140097944155080,
            outputs => outputs_140097944155080,
            outputs_full => outputs_full_140097944155080
        );
        
        core_inst_140097944155136: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944155136,
            fifo_full => fifo_full_140097944155136,
            outputs => outputs_140097944155136,
            outputs_full => outputs_full_140097944155136
        );
        
        core_inst_140097944155192: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944155192,
            fifo_full => fifo_full_140097944155192,
            outputs => outputs_140097944155192,
            outputs_full => outputs_full_140097944155192
        );
        
        core_inst_140097944155248: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944155248,
            fifo_full => fifo_full_140097944155248,
            outputs => outputs_140097944155248,
            outputs_full => outputs_full_140097944155248
        );
        
        core_inst_140097944155304: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944155304,
            fifo_full => fifo_full_140097944155304,
            outputs => outputs_140097944155304,
            outputs_full => outputs_full_140097944155304
        );
        
        core_inst_140097944155360: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944155360,
            fifo_full => fifo_full_140097944155360,
            outputs => outputs_140097944155360,
            outputs_full => outputs_full_140097944155360
        );
        
        core_inst_140097944155416: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944155416,
            fifo_full => fifo_full_140097944155416,
            outputs => outputs_140097944155416,
            outputs_full => outputs_full_140097944155416
        );
        
        core_inst_140097944155472: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944155472,
            fifo_full => fifo_full_140097944155472,
            outputs => outputs_140097944155472,
            outputs_full => outputs_full_140097944155472
        );
        
        core_inst_140097944155528: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944155528,
            fifo_full => fifo_full_140097944155528,
            outputs => outputs_140097944155528,
            outputs_full => outputs_full_140097944155528
        );
        
        core_inst_140097944155584: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944155584,
            fifo_full => fifo_full_140097944155584,
            outputs => outputs_140097944155584,
            outputs_full => outputs_full_140097944155584
        );
        
        core_inst_140097944155640: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944155640,
            fifo_full => fifo_full_140097944155640,
            outputs => outputs_140097944155640,
            outputs_full => outputs_full_140097944155640
        );
        
        core_inst_140097944155696: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944155696,
            fifo_full => fifo_full_140097944155696,
            outputs => outputs_140097944155696,
            outputs_full => outputs_full_140097944155696
        );
        
        core_inst_140097944155752: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944155752,
            fifo_full => fifo_full_140097944155752,
            outputs => outputs_140097944155752,
            outputs_full => outputs_full_140097944155752
        );
        
        core_inst_140097944155808: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944155808,
            fifo_full => fifo_full_140097944155808,
            outputs => outputs_140097944155808,
            outputs_full => outputs_full_140097944155808
        );
        
        core_inst_140097944155864: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944155864,
            fifo_full => fifo_full_140097944155864,
            outputs => outputs_140097944155864,
            outputs_full => outputs_full_140097944155864
        );
        
        core_inst_140097944155920: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944155920,
            fifo_full => fifo_full_140097944155920,
            outputs => outputs_140097944155920,
            outputs_full => outputs_full_140097944155920
        );
        
        core_inst_140097944155976: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944155976,
            fifo_full => fifo_full_140097944155976,
            outputs => outputs_140097944155976,
            outputs_full => outputs_full_140097944155976
        );
        
        core_inst_140097944156032: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944156032,
            fifo_full => fifo_full_140097944156032,
            outputs => outputs_140097944156032,
            outputs_full => outputs_full_140097944156032
        );
        
        core_inst_140097944156088: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944156088,
            fifo_full => fifo_full_140097944156088,
            outputs => outputs_140097944156088,
            outputs_full => outputs_full_140097944156088
        );
        
        core_inst_140097944156144: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944156144,
            fifo_full => fifo_full_140097944156144,
            outputs => outputs_140097944156144,
            outputs_full => outputs_full_140097944156144
        );
        
        core_inst_140097944156200: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944156200,
            fifo_full => fifo_full_140097944156200,
            outputs => outputs_140097944156200,
            outputs_full => outputs_full_140097944156200
        );
        
        core_inst_140097944156256: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944156256,
            fifo_full => fifo_full_140097944156256,
            outputs => outputs_140097944156256,
            outputs_full => outputs_full_140097944156256
        );
        
        core_inst_140097944156312: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944156312,
            fifo_full => fifo_full_140097944156312,
            outputs => outputs_140097944156312,
            outputs_full => outputs_full_140097944156312
        );
        
        core_inst_140097944156368: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944156368,
            fifo_full => fifo_full_140097944156368,
            outputs => outputs_140097944156368,
            outputs_full => outputs_full_140097944156368
        );
        
        core_inst_140097944156424: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944156424,
            fifo_full => fifo_full_140097944156424,
            outputs => outputs_140097944156424,
            outputs_full => outputs_full_140097944156424
        );
        
        core_inst_140097944156480: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944156480,
            fifo_full => fifo_full_140097944156480,
            outputs => outputs_140097944156480,
            outputs_full => outputs_full_140097944156480
        );
        
        core_inst_140097944156536: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944156536,
            fifo_full => fifo_full_140097944156536,
            outputs => outputs_140097944156536,
            outputs_full => outputs_full_140097944156536
        );
        
        core_inst_140097944156592: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944156592,
            fifo_full => fifo_full_140097944156592,
            outputs => outputs_140097944156592,
            outputs_full => outputs_full_140097944156592
        );
        
        core_inst_140097944156648: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944156648,
            fifo_full => fifo_full_140097944156648,
            outputs => outputs_140097944156648,
            outputs_full => outputs_full_140097944156648
        );
        
        core_inst_140097944156704: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944156704,
            fifo_full => fifo_full_140097944156704,
            outputs => outputs_140097944156704,
            outputs_full => outputs_full_140097944156704
        );
        
        core_inst_140097944156760: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944156760,
            fifo_full => fifo_full_140097944156760,
            outputs => outputs_140097944156760,
            outputs_full => outputs_full_140097944156760
        );
        
        core_inst_140097944156816: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944156816,
            fifo_full => fifo_full_140097944156816,
            outputs => outputs_140097944156816,
            outputs_full => outputs_full_140097944156816
        );
        
        core_inst_140097944156872: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944156872,
            fifo_full => fifo_full_140097944156872,
            outputs => outputs_140097944156872,
            outputs_full => outputs_full_140097944156872
        );
        
        core_inst_140097944156928: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944156928,
            fifo_full => fifo_full_140097944156928,
            outputs => outputs_140097944156928,
            outputs_full => outputs_full_140097944156928
        );
        
        core_inst_140097944156984: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944156984,
            fifo_full => fifo_full_140097944156984,
            outputs => outputs_140097944156984,
            outputs_full => outputs_full_140097944156984
        );
        
        core_inst_140097944157040: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944157040,
            fifo_full => fifo_full_140097944157040,
            outputs => outputs_140097944157040,
            outputs_full => outputs_full_140097944157040
        );
        
        core_inst_140097944157096: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944157096,
            fifo_full => fifo_full_140097944157096,
            outputs => outputs_140097944157096,
            outputs_full => outputs_full_140097944157096
        );
        
        core_inst_140097944157152: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944157152,
            fifo_full => fifo_full_140097944157152,
            outputs => outputs_140097944157152,
            outputs_full => outputs_full_140097944157152
        );
        
        core_inst_140097944157208: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944157208,
            fifo_full => fifo_full_140097944157208,
            outputs => outputs_140097944157208,
            outputs_full => outputs_full_140097944157208
        );
        
        core_inst_140097944157264: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944157264,
            fifo_full => fifo_full_140097944157264,
            outputs => outputs_140097944157264,
            outputs_full => outputs_full_140097944157264
        );
        
        core_inst_140097944157320: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944157320,
            fifo_full => fifo_full_140097944157320,
            outputs => outputs_140097944157320,
            outputs_full => outputs_full_140097944157320
        );
        
        core_inst_140097944157376: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944157376,
            fifo_full => fifo_full_140097944157376,
            outputs => outputs_140097944157376,
            outputs_full => outputs_full_140097944157376
        );
        
        core_inst_140097944157432: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944157432,
            fifo_full => fifo_full_140097944157432,
            outputs => outputs_140097944157432,
            outputs_full => outputs_full_140097944157432
        );
        
        core_inst_140097944157488: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944157488,
            fifo_full => fifo_full_140097944157488,
            outputs => outputs_140097944157488,
            outputs_full => outputs_full_140097944157488
        );
        
        core_inst_140097944157544: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944157544,
            fifo_full => fifo_full_140097944157544,
            outputs => outputs_140097944157544,
            outputs_full => outputs_full_140097944157544
        );
        
        core_inst_140097944157600: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944157600,
            fifo_full => fifo_full_140097944157600,
            outputs => outputs_140097944157600,
            outputs_full => outputs_full_140097944157600
        );
        
        core_inst_140097944157656: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944157656,
            fifo_full => fifo_full_140097944157656,
            outputs => outputs_140097944157656,
            outputs_full => outputs_full_140097944157656
        );
        
        core_inst_140097944157712: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944157712,
            fifo_full => fifo_full_140097944157712,
            outputs => outputs_140097944157712,
            outputs_full => outputs_full_140097944157712
        );
        
        core_inst_140097944157768: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944157768,
            fifo_full => fifo_full_140097944157768,
            outputs => outputs_140097944157768,
            outputs_full => outputs_full_140097944157768
        );
        
        core_inst_140097944157824: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944157824,
            fifo_full => fifo_full_140097944157824,
            outputs => outputs_140097944157824,
            outputs_full => outputs_full_140097944157824
        );
        
        core_inst_140097944157880: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944157880,
            fifo_full => fifo_full_140097944157880,
            outputs => outputs_140097944157880,
            outputs_full => outputs_full_140097944157880
        );
        
        core_inst_140097944157936: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944157936,
            fifo_full => fifo_full_140097944157936,
            outputs => outputs_140097944157936,
            outputs_full => outputs_full_140097944157936
        );
        
        core_inst_140097944157992: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944157992,
            fifo_full => fifo_full_140097944157992,
            outputs => outputs_140097944157992,
            outputs_full => outputs_full_140097944157992
        );
        
        core_inst_140097944158048: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944158048,
            fifo_full => fifo_full_140097944158048,
            outputs => outputs_140097944158048,
            outputs_full => outputs_full_140097944158048
        );
        
        core_inst_140097944158104: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944158104,
            fifo_full => fifo_full_140097944158104,
            outputs => outputs_140097944158104,
            outputs_full => outputs_full_140097944158104
        );
        
        core_inst_140097944158160: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944158160,
            fifo_full => fifo_full_140097944158160,
            outputs => outputs_140097944158160,
            outputs_full => outputs_full_140097944158160
        );
        
        core_inst_140097944166472: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944166472,
            fifo_full => fifo_full_140097944166472,
            outputs => outputs_140097944166472,
            outputs_full => outputs_full_140097944166472
        );
        
        core_inst_140097944166528: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944166528,
            fifo_full => fifo_full_140097944166528,
            outputs => outputs_140097944166528,
            outputs_full => outputs_full_140097944166528
        );
        
        core_inst_140097944166584: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944166584,
            fifo_full => fifo_full_140097944166584,
            outputs => outputs_140097944166584,
            outputs_full => outputs_full_140097944166584
        );
        
        core_inst_140097944166640: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944166640,
            fifo_full => fifo_full_140097944166640,
            outputs => outputs_140097944166640,
            outputs_full => outputs_full_140097944166640
        );
        
        core_inst_140097944166696: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944166696,
            fifo_full => fifo_full_140097944166696,
            outputs => outputs_140097944166696,
            outputs_full => outputs_full_140097944166696
        );
        
        core_inst_140097944166752: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944166752,
            fifo_full => fifo_full_140097944166752,
            outputs => outputs_140097944166752,
            outputs_full => outputs_full_140097944166752
        );
        
        core_inst_140097944166808: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944166808,
            fifo_full => fifo_full_140097944166808,
            outputs => outputs_140097944166808,
            outputs_full => outputs_full_140097944166808
        );
        
        core_inst_140097944166864: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944166864,
            fifo_full => fifo_full_140097944166864,
            outputs => outputs_140097944166864,
            outputs_full => outputs_full_140097944166864
        );
        
        core_inst_140097944166920: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944166920,
            fifo_full => fifo_full_140097944166920,
            outputs => outputs_140097944166920,
            outputs_full => outputs_full_140097944166920
        );
        
        core_inst_140097944166976: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944166976,
            fifo_full => fifo_full_140097944166976,
            outputs => outputs_140097944166976,
            outputs_full => outputs_full_140097944166976
        );
        
        core_inst_140097944167032: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944167032,
            fifo_full => fifo_full_140097944167032,
            outputs => outputs_140097944167032,
            outputs_full => outputs_full_140097944167032
        );
        
        core_inst_140097944167088: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944167088,
            fifo_full => fifo_full_140097944167088,
            outputs => outputs_140097944167088,
            outputs_full => outputs_full_140097944167088
        );
        
        core_inst_140097944167144: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944167144,
            fifo_full => fifo_full_140097944167144,
            outputs => outputs_140097944167144,
            outputs_full => outputs_full_140097944167144
        );
        
        core_inst_140097944167200: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944167200,
            fifo_full => fifo_full_140097944167200,
            outputs => outputs_140097944167200,
            outputs_full => outputs_full_140097944167200
        );
        
        core_inst_140097944167256: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944167256,
            fifo_full => fifo_full_140097944167256,
            outputs => outputs_140097944167256,
            outputs_full => outputs_full_140097944167256
        );
        
        core_inst_140097944167312: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944167312,
            fifo_full => fifo_full_140097944167312,
            outputs => outputs_140097944167312,
            outputs_full => outputs_full_140097944167312
        );
        
        core_inst_140097944167368: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944167368,
            fifo_full => fifo_full_140097944167368,
            outputs => outputs_140097944167368,
            outputs_full => outputs_full_140097944167368
        );
        
        core_inst_140097944167424: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944167424,
            fifo_full => fifo_full_140097944167424,
            outputs => outputs_140097944167424,
            outputs_full => outputs_full_140097944167424
        );
        
        core_inst_140097944167480: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944167480,
            fifo_full => fifo_full_140097944167480,
            outputs => outputs_140097944167480,
            outputs_full => outputs_full_140097944167480
        );
        
        core_inst_140097944167536: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944167536,
            fifo_full => fifo_full_140097944167536,
            outputs => outputs_140097944167536,
            outputs_full => outputs_full_140097944167536
        );
        
        core_inst_140097944167592: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944167592,
            fifo_full => fifo_full_140097944167592,
            outputs => outputs_140097944167592,
            outputs_full => outputs_full_140097944167592
        );
        
        core_inst_140097944167648: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944167648,
            fifo_full => fifo_full_140097944167648,
            outputs => outputs_140097944167648,
            outputs_full => outputs_full_140097944167648
        );
        
        core_inst_140097944167704: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944167704,
            fifo_full => fifo_full_140097944167704,
            outputs => outputs_140097944167704,
            outputs_full => outputs_full_140097944167704
        );
        
        core_inst_140097944167760: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944167760,
            fifo_full => fifo_full_140097944167760,
            outputs => outputs_140097944167760,
            outputs_full => outputs_full_140097944167760
        );
        
        core_inst_140097944167816: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944167816,
            fifo_full => fifo_full_140097944167816,
            outputs => outputs_140097944167816,
            outputs_full => outputs_full_140097944167816
        );
        
        core_inst_140097944167872: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944167872,
            fifo_full => fifo_full_140097944167872,
            outputs => outputs_140097944167872,
            outputs_full => outputs_full_140097944167872
        );
        
        core_inst_140097944167928: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944167928,
            fifo_full => fifo_full_140097944167928,
            outputs => outputs_140097944167928,
            outputs_full => outputs_full_140097944167928
        );
        
        core_inst_140097944167984: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944167984,
            fifo_full => fifo_full_140097944167984,
            outputs => outputs_140097944167984,
            outputs_full => outputs_full_140097944167984
        );
        
        core_inst_140097944168040: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944168040,
            fifo_full => fifo_full_140097944168040,
            outputs => outputs_140097944168040,
            outputs_full => outputs_full_140097944168040
        );
        
        core_inst_140097944168096: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944168096,
            fifo_full => fifo_full_140097944168096,
            outputs => outputs_140097944168096,
            outputs_full => outputs_full_140097944168096
        );
        
        core_inst_140097944168152: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944168152,
            fifo_full => fifo_full_140097944168152,
            outputs => outputs_140097944168152,
            outputs_full => outputs_full_140097944168152
        );
        
        core_inst_140097944168208: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944168208,
            fifo_full => fifo_full_140097944168208,
            outputs => outputs_140097944168208,
            outputs_full => outputs_full_140097944168208
        );
        
        core_inst_140097944168264: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944168264,
            fifo_full => fifo_full_140097944168264,
            outputs => outputs_140097944168264,
            outputs_full => outputs_full_140097944168264
        );
        
        core_inst_140097944168320: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944168320,
            fifo_full => fifo_full_140097944168320,
            outputs => outputs_140097944168320,
            outputs_full => outputs_full_140097944168320
        );
        
        core_inst_140097944168376: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944168376,
            fifo_full => fifo_full_140097944168376,
            outputs => outputs_140097944168376,
            outputs_full => outputs_full_140097944168376
        );
        
        core_inst_140097944168432: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944168432,
            fifo_full => fifo_full_140097944168432,
            outputs => outputs_140097944168432,
            outputs_full => outputs_full_140097944168432
        );
        
        core_inst_140097944168488: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944168488,
            fifo_full => fifo_full_140097944168488,
            outputs => outputs_140097944168488,
            outputs_full => outputs_full_140097944168488
        );
        
        core_inst_140097944168544: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944168544,
            fifo_full => fifo_full_140097944168544,
            outputs => outputs_140097944168544,
            outputs_full => outputs_full_140097944168544
        );
        
        core_inst_140097944168600: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944168600,
            fifo_full => fifo_full_140097944168600,
            outputs => outputs_140097944168600,
            outputs_full => outputs_full_140097944168600
        );
        
        core_inst_140097944168656: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944168656,
            fifo_full => fifo_full_140097944168656,
            outputs => outputs_140097944168656,
            outputs_full => outputs_full_140097944168656
        );
        
        core_inst_140097944168712: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944168712,
            fifo_full => fifo_full_140097944168712,
            outputs => outputs_140097944168712,
            outputs_full => outputs_full_140097944168712
        );
        
        core_inst_140097944168768: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944168768,
            fifo_full => fifo_full_140097944168768,
            outputs => outputs_140097944168768,
            outputs_full => outputs_full_140097944168768
        );
        
        core_inst_140097944168824: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944168824,
            fifo_full => fifo_full_140097944168824,
            outputs => outputs_140097944168824,
            outputs_full => outputs_full_140097944168824
        );
        
        core_inst_140097944168880: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944168880,
            fifo_full => fifo_full_140097944168880,
            outputs => outputs_140097944168880,
            outputs_full => outputs_full_140097944168880
        );
        
        core_inst_140097944168936: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944168936,
            fifo_full => fifo_full_140097944168936,
            outputs => outputs_140097944168936,
            outputs_full => outputs_full_140097944168936
        );
        
        core_inst_140097944168992: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944168992,
            fifo_full => fifo_full_140097944168992,
            outputs => outputs_140097944168992,
            outputs_full => outputs_full_140097944168992
        );
        
        core_inst_140097944169048: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944169048,
            fifo_full => fifo_full_140097944169048,
            outputs => outputs_140097944169048,
            outputs_full => outputs_full_140097944169048
        );
        
        core_inst_140097944169104: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944169104,
            fifo_full => fifo_full_140097944169104,
            outputs => outputs_140097944169104,
            outputs_full => outputs_full_140097944169104
        );
        
        core_inst_140097944169160: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944169160,
            fifo_full => fifo_full_140097944169160,
            outputs => outputs_140097944169160,
            outputs_full => outputs_full_140097944169160
        );
        
        core_inst_140097944169216: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944169216,
            fifo_full => fifo_full_140097944169216,
            outputs => outputs_140097944169216,
            outputs_full => outputs_full_140097944169216
        );
        
        core_inst_140097944169272: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944169272,
            fifo_full => fifo_full_140097944169272,
            outputs => outputs_140097944169272,
            outputs_full => outputs_full_140097944169272
        );
        
        core_inst_140097944169328: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944169328,
            fifo_full => fifo_full_140097944169328,
            outputs => outputs_140097944169328,
            outputs_full => outputs_full_140097944169328
        );
        
        core_inst_140097944169384: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944169384,
            fifo_full => fifo_full_140097944169384,
            outputs => outputs_140097944169384,
            outputs_full => outputs_full_140097944169384
        );
        
        core_inst_140097944169440: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944169440,
            fifo_full => fifo_full_140097944169440,
            outputs => outputs_140097944169440,
            outputs_full => outputs_full_140097944169440
        );
        
        core_inst_140097944169496: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944169496,
            fifo_full => fifo_full_140097944169496,
            outputs => outputs_140097944169496,
            outputs_full => outputs_full_140097944169496
        );
        
        core_inst_140097944169552: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944169552,
            fifo_full => fifo_full_140097944169552,
            outputs => outputs_140097944169552,
            outputs_full => outputs_full_140097944169552
        );
        
        core_inst_140097944169608: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944169608,
            fifo_full => fifo_full_140097944169608,
            outputs => outputs_140097944169608,
            outputs_full => outputs_full_140097944169608
        );
        
        core_inst_140097944169664: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944169664,
            fifo_full => fifo_full_140097944169664,
            outputs => outputs_140097944169664,
            outputs_full => outputs_full_140097944169664
        );
        
        core_inst_140097944169720: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944169720,
            fifo_full => fifo_full_140097944169720,
            outputs => outputs_140097944169720,
            outputs_full => outputs_full_140097944169720
        );
        
        core_inst_140097944169776: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944169776,
            fifo_full => fifo_full_140097944169776,
            outputs => outputs_140097944169776,
            outputs_full => outputs_full_140097944169776
        );
        
        core_inst_140097944169832: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944169832,
            fifo_full => fifo_full_140097944169832,
            outputs => outputs_140097944169832,
            outputs_full => outputs_full_140097944169832
        );
        
        core_inst_140097944169888: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944169888,
            fifo_full => fifo_full_140097944169888,
            outputs => outputs_140097944169888,
            outputs_full => outputs_full_140097944169888
        );
        
        core_inst_140097944169944: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944169944,
            fifo_full => fifo_full_140097944169944,
            outputs => outputs_140097944169944,
            outputs_full => outputs_full_140097944169944
        );
        
        core_inst_140097944170000: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944170000,
            fifo_full => fifo_full_140097944170000,
            outputs => outputs_140097944170000,
            outputs_full => outputs_full_140097944170000
        );
        
        core_inst_140097944170056: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944170056,
            fifo_full => fifo_full_140097944170056,
            outputs => outputs_140097944170056,
            outputs_full => outputs_full_140097944170056
        );
        
        core_inst_140097944170112: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944170112,
            fifo_full => fifo_full_140097944170112,
            outputs => outputs_140097944170112,
            outputs_full => outputs_full_140097944170112
        );
        
        core_inst_140097944170168: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944170168,
            fifo_full => fifo_full_140097944170168,
            outputs => outputs_140097944170168,
            outputs_full => outputs_full_140097944170168
        );
        
        core_inst_140097944170224: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944170224,
            fifo_full => fifo_full_140097944170224,
            outputs => outputs_140097944170224,
            outputs_full => outputs_full_140097944170224
        );
        
        core_inst_140097944170280: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944170280,
            fifo_full => fifo_full_140097944170280,
            outputs => outputs_140097944170280,
            outputs_full => outputs_full_140097944170280
        );
        
        core_inst_140097944170336: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944170336,
            fifo_full => fifo_full_140097944170336,
            outputs => outputs_140097944170336,
            outputs_full => outputs_full_140097944170336
        );
        
        core_inst_140097944170392: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944170392,
            fifo_full => fifo_full_140097944170392,
            outputs => outputs_140097944170392,
            outputs_full => outputs_full_140097944170392
        );
        
        core_inst_140097944170448: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097944170448,
            fifo_full => fifo_full_140097944170448,
            outputs => outputs_140097944170448,
            outputs_full => outputs_full_140097944170448
        );
        
        core_inst_140097941516360: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941516360,
            fifo_full => fifo_full_140097941516360,
            outputs => outputs_140097941516360,
            outputs_full => outputs_full_140097941516360
        );
        
        core_inst_140097941516416: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941516416,
            fifo_full => fifo_full_140097941516416,
            outputs => outputs_140097941516416,
            outputs_full => outputs_full_140097941516416
        );
        
        core_inst_140097941516472: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941516472,
            fifo_full => fifo_full_140097941516472,
            outputs => outputs_140097941516472,
            outputs_full => outputs_full_140097941516472
        );
        
        core_inst_140097941516528: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941516528,
            fifo_full => fifo_full_140097941516528,
            outputs => outputs_140097941516528,
            outputs_full => outputs_full_140097941516528
        );
        
        core_inst_140097941516584: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941516584,
            fifo_full => fifo_full_140097941516584,
            outputs => outputs_140097941516584,
            outputs_full => outputs_full_140097941516584
        );
        
        core_inst_140097941516640: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941516640,
            fifo_full => fifo_full_140097941516640,
            outputs => outputs_140097941516640,
            outputs_full => outputs_full_140097941516640
        );
        
        core_inst_140097941516696: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941516696,
            fifo_full => fifo_full_140097941516696,
            outputs => outputs_140097941516696,
            outputs_full => outputs_full_140097941516696
        );
        
        core_inst_140097941516752: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941516752,
            fifo_full => fifo_full_140097941516752,
            outputs => outputs_140097941516752,
            outputs_full => outputs_full_140097941516752
        );
        
        core_inst_140097941516808: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941516808,
            fifo_full => fifo_full_140097941516808,
            outputs => outputs_140097941516808,
            outputs_full => outputs_full_140097941516808
        );
        
        core_inst_140097941516864: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941516864,
            fifo_full => fifo_full_140097941516864,
            outputs => outputs_140097941516864,
            outputs_full => outputs_full_140097941516864
        );
        
        core_inst_140097941516920: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941516920,
            fifo_full => fifo_full_140097941516920,
            outputs => outputs_140097941516920,
            outputs_full => outputs_full_140097941516920
        );
        
        core_inst_140097941516976: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941516976,
            fifo_full => fifo_full_140097941516976,
            outputs => outputs_140097941516976,
            outputs_full => outputs_full_140097941516976
        );
        
        core_inst_140097941517032: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941517032,
            fifo_full => fifo_full_140097941517032,
            outputs => outputs_140097941517032,
            outputs_full => outputs_full_140097941517032
        );
        
        core_inst_140097941517088: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941517088,
            fifo_full => fifo_full_140097941517088,
            outputs => outputs_140097941517088,
            outputs_full => outputs_full_140097941517088
        );
        
        core_inst_140097941517144: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941517144,
            fifo_full => fifo_full_140097941517144,
            outputs => outputs_140097941517144,
            outputs_full => outputs_full_140097941517144
        );
        
        core_inst_140097941517200: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941517200,
            fifo_full => fifo_full_140097941517200,
            outputs => outputs_140097941517200,
            outputs_full => outputs_full_140097941517200
        );
        
        core_inst_140097941517256: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941517256,
            fifo_full => fifo_full_140097941517256,
            outputs => outputs_140097941517256,
            outputs_full => outputs_full_140097941517256
        );
        
        core_inst_140097941517312: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941517312,
            fifo_full => fifo_full_140097941517312,
            outputs => outputs_140097941517312,
            outputs_full => outputs_full_140097941517312
        );
        
        core_inst_140097941517368: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941517368,
            fifo_full => fifo_full_140097941517368,
            outputs => outputs_140097941517368,
            outputs_full => outputs_full_140097941517368
        );
        
        core_inst_140097941517424: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941517424,
            fifo_full => fifo_full_140097941517424,
            outputs => outputs_140097941517424,
            outputs_full => outputs_full_140097941517424
        );
        
        core_inst_140097941517480: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941517480,
            fifo_full => fifo_full_140097941517480,
            outputs => outputs_140097941517480,
            outputs_full => outputs_full_140097941517480
        );
        
        core_inst_140097941517536: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941517536,
            fifo_full => fifo_full_140097941517536,
            outputs => outputs_140097941517536,
            outputs_full => outputs_full_140097941517536
        );
        
        core_inst_140097941517592: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941517592,
            fifo_full => fifo_full_140097941517592,
            outputs => outputs_140097941517592,
            outputs_full => outputs_full_140097941517592
        );
        
        core_inst_140097941517648: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941517648,
            fifo_full => fifo_full_140097941517648,
            outputs => outputs_140097941517648,
            outputs_full => outputs_full_140097941517648
        );
        
        core_inst_140097941517704: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941517704,
            fifo_full => fifo_full_140097941517704,
            outputs => outputs_140097941517704,
            outputs_full => outputs_full_140097941517704
        );
        
        core_inst_140097941517760: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941517760,
            fifo_full => fifo_full_140097941517760,
            outputs => outputs_140097941517760,
            outputs_full => outputs_full_140097941517760
        );
        
        core_inst_140097941517816: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941517816,
            fifo_full => fifo_full_140097941517816,
            outputs => outputs_140097941517816,
            outputs_full => outputs_full_140097941517816
        );
        
        core_inst_140097941517872: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941517872,
            fifo_full => fifo_full_140097941517872,
            outputs => outputs_140097941517872,
            outputs_full => outputs_full_140097941517872
        );
        
        core_inst_140097941517928: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941517928,
            fifo_full => fifo_full_140097941517928,
            outputs => outputs_140097941517928,
            outputs_full => outputs_full_140097941517928
        );
        
        core_inst_140097941517984: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941517984,
            fifo_full => fifo_full_140097941517984,
            outputs => outputs_140097941517984,
            outputs_full => outputs_full_140097941517984
        );
        
        core_inst_140097941518040: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941518040,
            fifo_full => fifo_full_140097941518040,
            outputs => outputs_140097941518040,
            outputs_full => outputs_full_140097941518040
        );
        
        core_inst_140097941518096: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941518096,
            fifo_full => fifo_full_140097941518096,
            outputs => outputs_140097941518096,
            outputs_full => outputs_full_140097941518096
        );
        
        core_inst_140097941518152: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941518152,
            fifo_full => fifo_full_140097941518152,
            outputs => outputs_140097941518152,
            outputs_full => outputs_full_140097941518152
        );
        
        core_inst_140097941518208: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941518208,
            fifo_full => fifo_full_140097941518208,
            outputs => outputs_140097941518208,
            outputs_full => outputs_full_140097941518208
        );
        
        core_inst_140097941518264: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941518264,
            fifo_full => fifo_full_140097941518264,
            outputs => outputs_140097941518264,
            outputs_full => outputs_full_140097941518264
        );
        
        core_inst_140097941518320: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941518320,
            fifo_full => fifo_full_140097941518320,
            outputs => outputs_140097941518320,
            outputs_full => outputs_full_140097941518320
        );
        
        core_inst_140097941518376: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941518376,
            fifo_full => fifo_full_140097941518376,
            outputs => outputs_140097941518376,
            outputs_full => outputs_full_140097941518376
        );
        
        core_inst_140097941518432: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941518432,
            fifo_full => fifo_full_140097941518432,
            outputs => outputs_140097941518432,
            outputs_full => outputs_full_140097941518432
        );
        
        core_inst_140097941518488: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941518488,
            fifo_full => fifo_full_140097941518488,
            outputs => outputs_140097941518488,
            outputs_full => outputs_full_140097941518488
        );
        
        core_inst_140097941518544: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941518544,
            fifo_full => fifo_full_140097941518544,
            outputs => outputs_140097941518544,
            outputs_full => outputs_full_140097941518544
        );
        
        core_inst_140097941518600: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941518600,
            fifo_full => fifo_full_140097941518600,
            outputs => outputs_140097941518600,
            outputs_full => outputs_full_140097941518600
        );
        
        core_inst_140097941518656: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941518656,
            fifo_full => fifo_full_140097941518656,
            outputs => outputs_140097941518656,
            outputs_full => outputs_full_140097941518656
        );
        
        core_inst_140097941518712: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941518712,
            fifo_full => fifo_full_140097941518712,
            outputs => outputs_140097941518712,
            outputs_full => outputs_full_140097941518712
        );
        
        core_inst_140097941518768: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941518768,
            fifo_full => fifo_full_140097941518768,
            outputs => outputs_140097941518768,
            outputs_full => outputs_full_140097941518768
        );
        
        core_inst_140097941518824: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941518824,
            fifo_full => fifo_full_140097941518824,
            outputs => outputs_140097941518824,
            outputs_full => outputs_full_140097941518824
        );
        
        core_inst_140097941518880: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941518880,
            fifo_full => fifo_full_140097941518880,
            outputs => outputs_140097941518880,
            outputs_full => outputs_full_140097941518880
        );
        
        core_inst_140097941518936: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941518936,
            fifo_full => fifo_full_140097941518936,
            outputs => outputs_140097941518936,
            outputs_full => outputs_full_140097941518936
        );
        
        core_inst_140097941518992: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941518992,
            fifo_full => fifo_full_140097941518992,
            outputs => outputs_140097941518992,
            outputs_full => outputs_full_140097941518992
        );
        
        core_inst_140097941519048: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941519048,
            fifo_full => fifo_full_140097941519048,
            outputs => outputs_140097941519048,
            outputs_full => outputs_full_140097941519048
        );
        
        core_inst_140097941519104: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941519104,
            fifo_full => fifo_full_140097941519104,
            outputs => outputs_140097941519104,
            outputs_full => outputs_full_140097941519104
        );
        
        core_inst_140097941519160: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941519160,
            fifo_full => fifo_full_140097941519160,
            outputs => outputs_140097941519160,
            outputs_full => outputs_full_140097941519160
        );
        
        core_inst_140097941519216: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941519216,
            fifo_full => fifo_full_140097941519216,
            outputs => outputs_140097941519216,
            outputs_full => outputs_full_140097941519216
        );
        
        core_inst_140097941519272: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941519272,
            fifo_full => fifo_full_140097941519272,
            outputs => outputs_140097941519272,
            outputs_full => outputs_full_140097941519272
        );
        
        core_inst_140097941519328: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941519328,
            fifo_full => fifo_full_140097941519328,
            outputs => outputs_140097941519328,
            outputs_full => outputs_full_140097941519328
        );
        
        core_inst_140097941519384: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941519384,
            fifo_full => fifo_full_140097941519384,
            outputs => outputs_140097941519384,
            outputs_full => outputs_full_140097941519384
        );
        
        core_inst_140097941519440: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941519440,
            fifo_full => fifo_full_140097941519440,
            outputs => outputs_140097941519440,
            outputs_full => outputs_full_140097941519440
        );
        
        core_inst_140097941519496: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941519496,
            fifo_full => fifo_full_140097941519496,
            outputs => outputs_140097941519496,
            outputs_full => outputs_full_140097941519496
        );
        
        core_inst_140097941519552: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941519552,
            fifo_full => fifo_full_140097941519552,
            outputs => outputs_140097941519552,
            outputs_full => outputs_full_140097941519552
        );
        
        core_inst_140097941519608: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941519608,
            fifo_full => fifo_full_140097941519608,
            outputs => outputs_140097941519608,
            outputs_full => outputs_full_140097941519608
        );
        
        core_inst_140097941519664: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941519664,
            fifo_full => fifo_full_140097941519664,
            outputs => outputs_140097941519664,
            outputs_full => outputs_full_140097941519664
        );
        
        core_inst_140097941519720: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941519720,
            fifo_full => fifo_full_140097941519720,
            outputs => outputs_140097941519720,
            outputs_full => outputs_full_140097941519720
        );
        
        core_inst_140097941519776: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941519776,
            fifo_full => fifo_full_140097941519776,
            outputs => outputs_140097941519776,
            outputs_full => outputs_full_140097941519776
        );
        
        core_inst_140097941519832: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941519832,
            fifo_full => fifo_full_140097941519832,
            outputs => outputs_140097941519832,
            outputs_full => outputs_full_140097941519832
        );
        
        core_inst_140097941519888: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941519888,
            fifo_full => fifo_full_140097941519888,
            outputs => outputs_140097941519888,
            outputs_full => outputs_full_140097941519888
        );
        
        core_inst_140097941519944: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941519944,
            fifo_full => fifo_full_140097941519944,
            outputs => outputs_140097941519944,
            outputs_full => outputs_full_140097941519944
        );
        
        core_inst_140097941520000: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941520000,
            fifo_full => fifo_full_140097941520000,
            outputs => outputs_140097941520000,
            outputs_full => outputs_full_140097941520000
        );
        
        core_inst_140097941520056: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941520056,
            fifo_full => fifo_full_140097941520056,
            outputs => outputs_140097941520056,
            outputs_full => outputs_full_140097941520056
        );
        
        core_inst_140097941520112: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941520112,
            fifo_full => fifo_full_140097941520112,
            outputs => outputs_140097941520112,
            outputs_full => outputs_full_140097941520112
        );
        
        core_inst_140097941520168: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941520168,
            fifo_full => fifo_full_140097941520168,
            outputs => outputs_140097941520168,
            outputs_full => outputs_full_140097941520168
        );
        
        core_inst_140097941520224: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941520224,
            fifo_full => fifo_full_140097941520224,
            outputs => outputs_140097941520224,
            outputs_full => outputs_full_140097941520224
        );
        
        core_inst_140097941520280: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941520280,
            fifo_full => fifo_full_140097941520280,
            outputs => outputs_140097941520280,
            outputs_full => outputs_full_140097941520280
        );
        
        core_inst_140097941520336: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941520336,
            fifo_full => fifo_full_140097941520336,
            outputs => outputs_140097941520336,
            outputs_full => outputs_full_140097941520336
        );
        
        core_inst_140097941528648: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941528648,
            fifo_full => fifo_full_140097941528648,
            outputs => outputs_140097941528648,
            outputs_full => outputs_full_140097941528648
        );
        
        core_inst_140097941528704: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941528704,
            fifo_full => fifo_full_140097941528704,
            outputs => outputs_140097941528704,
            outputs_full => outputs_full_140097941528704
        );
        
        core_inst_140097941528760: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941528760,
            fifo_full => fifo_full_140097941528760,
            outputs => outputs_140097941528760,
            outputs_full => outputs_full_140097941528760
        );
        
        core_inst_140097941528816: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941528816,
            fifo_full => fifo_full_140097941528816,
            outputs => outputs_140097941528816,
            outputs_full => outputs_full_140097941528816
        );
        
        core_inst_140097941528872: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941528872,
            fifo_full => fifo_full_140097941528872,
            outputs => outputs_140097941528872,
            outputs_full => outputs_full_140097941528872
        );
        
        core_inst_140097941528928: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941528928,
            fifo_full => fifo_full_140097941528928,
            outputs => outputs_140097941528928,
            outputs_full => outputs_full_140097941528928
        );
        
        core_inst_140097941528984: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941528984,
            fifo_full => fifo_full_140097941528984,
            outputs => outputs_140097941528984,
            outputs_full => outputs_full_140097941528984
        );
        
        core_inst_140097941529040: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941529040,
            fifo_full => fifo_full_140097941529040,
            outputs => outputs_140097941529040,
            outputs_full => outputs_full_140097941529040
        );
        
        core_inst_140097941529096: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941529096,
            fifo_full => fifo_full_140097941529096,
            outputs => outputs_140097941529096,
            outputs_full => outputs_full_140097941529096
        );
        
        core_inst_140097941529152: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941529152,
            fifo_full => fifo_full_140097941529152,
            outputs => outputs_140097941529152,
            outputs_full => outputs_full_140097941529152
        );
        
        core_inst_140097941529208: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941529208,
            fifo_full => fifo_full_140097941529208,
            outputs => outputs_140097941529208,
            outputs_full => outputs_full_140097941529208
        );
        
        core_inst_140097941529264: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941529264,
            fifo_full => fifo_full_140097941529264,
            outputs => outputs_140097941529264,
            outputs_full => outputs_full_140097941529264
        );
        
        core_inst_140097941529320: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941529320,
            fifo_full => fifo_full_140097941529320,
            outputs => outputs_140097941529320,
            outputs_full => outputs_full_140097941529320
        );
        
        core_inst_140097941529376: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941529376,
            fifo_full => fifo_full_140097941529376,
            outputs => outputs_140097941529376,
            outputs_full => outputs_full_140097941529376
        );
        
        core_inst_140097941529432: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941529432,
            fifo_full => fifo_full_140097941529432,
            outputs => outputs_140097941529432,
            outputs_full => outputs_full_140097941529432
        );
        
        core_inst_140097941529488: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941529488,
            fifo_full => fifo_full_140097941529488,
            outputs => outputs_140097941529488,
            outputs_full => outputs_full_140097941529488
        );
        
        core_inst_140097941529544: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941529544,
            fifo_full => fifo_full_140097941529544,
            outputs => outputs_140097941529544,
            outputs_full => outputs_full_140097941529544
        );
        
        core_inst_140097941529600: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941529600,
            fifo_full => fifo_full_140097941529600,
            outputs => outputs_140097941529600,
            outputs_full => outputs_full_140097941529600
        );
        
        core_inst_140097941529656: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941529656,
            fifo_full => fifo_full_140097941529656,
            outputs => outputs_140097941529656,
            outputs_full => outputs_full_140097941529656
        );
        
        core_inst_140097941529712: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941529712,
            fifo_full => fifo_full_140097941529712,
            outputs => outputs_140097941529712,
            outputs_full => outputs_full_140097941529712
        );
        
        core_inst_140097941529768: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941529768,
            fifo_full => fifo_full_140097941529768,
            outputs => outputs_140097941529768,
            outputs_full => outputs_full_140097941529768
        );
        
        core_inst_140097941529824: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941529824,
            fifo_full => fifo_full_140097941529824,
            outputs => outputs_140097941529824,
            outputs_full => outputs_full_140097941529824
        );
        
        core_inst_140097941529880: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941529880,
            fifo_full => fifo_full_140097941529880,
            outputs => outputs_140097941529880,
            outputs_full => outputs_full_140097941529880
        );
        
        core_inst_140097941529936: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941529936,
            fifo_full => fifo_full_140097941529936,
            outputs => outputs_140097941529936,
            outputs_full => outputs_full_140097941529936
        );
        
        core_inst_140097941529992: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941529992,
            fifo_full => fifo_full_140097941529992,
            outputs => outputs_140097941529992,
            outputs_full => outputs_full_140097941529992
        );
        
        core_inst_140097941530048: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941530048,
            fifo_full => fifo_full_140097941530048,
            outputs => outputs_140097941530048,
            outputs_full => outputs_full_140097941530048
        );
        
        core_inst_140097941530104: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941530104,
            fifo_full => fifo_full_140097941530104,
            outputs => outputs_140097941530104,
            outputs_full => outputs_full_140097941530104
        );
        
        core_inst_140097941530160: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941530160,
            fifo_full => fifo_full_140097941530160,
            outputs => outputs_140097941530160,
            outputs_full => outputs_full_140097941530160
        );
        
        core_inst_140097941530216: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941530216,
            fifo_full => fifo_full_140097941530216,
            outputs => outputs_140097941530216,
            outputs_full => outputs_full_140097941530216
        );
        
        core_inst_140097941530272: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941530272,
            fifo_full => fifo_full_140097941530272,
            outputs => outputs_140097941530272,
            outputs_full => outputs_full_140097941530272
        );
        
        core_inst_140097941530328: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941530328,
            fifo_full => fifo_full_140097941530328,
            outputs => outputs_140097941530328,
            outputs_full => outputs_full_140097941530328
        );
        
        core_inst_140097941530384: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941530384,
            fifo_full => fifo_full_140097941530384,
            outputs => outputs_140097941530384,
            outputs_full => outputs_full_140097941530384
        );
        
        core_inst_140097941530440: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941530440,
            fifo_full => fifo_full_140097941530440,
            outputs => outputs_140097941530440,
            outputs_full => outputs_full_140097941530440
        );
        
        core_inst_140097941530496: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941530496,
            fifo_full => fifo_full_140097941530496,
            outputs => outputs_140097941530496,
            outputs_full => outputs_full_140097941530496
        );
        
        core_inst_140097941530552: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941530552,
            fifo_full => fifo_full_140097941530552,
            outputs => outputs_140097941530552,
            outputs_full => outputs_full_140097941530552
        );
        
        core_inst_140097941530608: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941530608,
            fifo_full => fifo_full_140097941530608,
            outputs => outputs_140097941530608,
            outputs_full => outputs_full_140097941530608
        );
        
        core_inst_140097941530664: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941530664,
            fifo_full => fifo_full_140097941530664,
            outputs => outputs_140097941530664,
            outputs_full => outputs_full_140097941530664
        );
        
        core_inst_140097941530720: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941530720,
            fifo_full => fifo_full_140097941530720,
            outputs => outputs_140097941530720,
            outputs_full => outputs_full_140097941530720
        );
        
        core_inst_140097941530776: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941530776,
            fifo_full => fifo_full_140097941530776,
            outputs => outputs_140097941530776,
            outputs_full => outputs_full_140097941530776
        );
        
        core_inst_140097941530832: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941530832,
            fifo_full => fifo_full_140097941530832,
            outputs => outputs_140097941530832,
            outputs_full => outputs_full_140097941530832
        );
        
        core_inst_140097941530888: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941530888,
            fifo_full => fifo_full_140097941530888,
            outputs => outputs_140097941530888,
            outputs_full => outputs_full_140097941530888
        );
        
        core_inst_140097941530944: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941530944,
            fifo_full => fifo_full_140097941530944,
            outputs => outputs_140097941530944,
            outputs_full => outputs_full_140097941530944
        );
        
        core_inst_140097941531000: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941531000,
            fifo_full => fifo_full_140097941531000,
            outputs => outputs_140097941531000,
            outputs_full => outputs_full_140097941531000
        );
        
        core_inst_140097941531056: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941531056,
            fifo_full => fifo_full_140097941531056,
            outputs => outputs_140097941531056,
            outputs_full => outputs_full_140097941531056
        );
        
        core_inst_140097941531112: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941531112,
            fifo_full => fifo_full_140097941531112,
            outputs => outputs_140097941531112,
            outputs_full => outputs_full_140097941531112
        );
        
        core_inst_140097941531168: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941531168,
            fifo_full => fifo_full_140097941531168,
            outputs => outputs_140097941531168,
            outputs_full => outputs_full_140097941531168
        );
        
        core_inst_140097941531224: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941531224,
            fifo_full => fifo_full_140097941531224,
            outputs => outputs_140097941531224,
            outputs_full => outputs_full_140097941531224
        );
        
        core_inst_140097941531280: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941531280,
            fifo_full => fifo_full_140097941531280,
            outputs => outputs_140097941531280,
            outputs_full => outputs_full_140097941531280
        );
        
        core_inst_140097941531336: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941531336,
            fifo_full => fifo_full_140097941531336,
            outputs => outputs_140097941531336,
            outputs_full => outputs_full_140097941531336
        );
        
        core_inst_140097941531392: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941531392,
            fifo_full => fifo_full_140097941531392,
            outputs => outputs_140097941531392,
            outputs_full => outputs_full_140097941531392
        );
        
        core_inst_140097941531448: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941531448,
            fifo_full => fifo_full_140097941531448,
            outputs => outputs_140097941531448,
            outputs_full => outputs_full_140097941531448
        );
        
        core_inst_140097941531504: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941531504,
            fifo_full => fifo_full_140097941531504,
            outputs => outputs_140097941531504,
            outputs_full => outputs_full_140097941531504
        );
        
        core_inst_140097941531560: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941531560,
            fifo_full => fifo_full_140097941531560,
            outputs => outputs_140097941531560,
            outputs_full => outputs_full_140097941531560
        );
        
        core_inst_140097941531616: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941531616,
            fifo_full => fifo_full_140097941531616,
            outputs => outputs_140097941531616,
            outputs_full => outputs_full_140097941531616
        );
        
        core_inst_140097941531672: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941531672,
            fifo_full => fifo_full_140097941531672,
            outputs => outputs_140097941531672,
            outputs_full => outputs_full_140097941531672
        );
        
        core_inst_140097941531728: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941531728,
            fifo_full => fifo_full_140097941531728,
            outputs => outputs_140097941531728,
            outputs_full => outputs_full_140097941531728
        );
        
        core_inst_140097941531784: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941531784,
            fifo_full => fifo_full_140097941531784,
            outputs => outputs_140097941531784,
            outputs_full => outputs_full_140097941531784
        );
        
        core_inst_140097941531840: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941531840,
            fifo_full => fifo_full_140097941531840,
            outputs => outputs_140097941531840,
            outputs_full => outputs_full_140097941531840
        );
        
        core_inst_140097941531896: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941531896,
            fifo_full => fifo_full_140097941531896,
            outputs => outputs_140097941531896,
            outputs_full => outputs_full_140097941531896
        );
        
        core_inst_140097941531952: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941531952,
            fifo_full => fifo_full_140097941531952,
            outputs => outputs_140097941531952,
            outputs_full => outputs_full_140097941531952
        );
        
        core_inst_140097941532008: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941532008,
            fifo_full => fifo_full_140097941532008,
            outputs => outputs_140097941532008,
            outputs_full => outputs_full_140097941532008
        );
        
        core_inst_140097941532064: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941532064,
            fifo_full => fifo_full_140097941532064,
            outputs => outputs_140097941532064,
            outputs_full => outputs_full_140097941532064
        );
        
        core_inst_140097941532120: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941532120,
            fifo_full => fifo_full_140097941532120,
            outputs => outputs_140097941532120,
            outputs_full => outputs_full_140097941532120
        );
        
        core_inst_140097941532176: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941532176,
            fifo_full => fifo_full_140097941532176,
            outputs => outputs_140097941532176,
            outputs_full => outputs_full_140097941532176
        );
        
        core_inst_140097941532232: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941532232,
            fifo_full => fifo_full_140097941532232,
            outputs => outputs_140097941532232,
            outputs_full => outputs_full_140097941532232
        );
        
        core_inst_140097941532288: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941532288,
            fifo_full => fifo_full_140097941532288,
            outputs => outputs_140097941532288,
            outputs_full => outputs_full_140097941532288
        );
        
        core_inst_140097941532344: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941532344,
            fifo_full => fifo_full_140097941532344,
            outputs => outputs_140097941532344,
            outputs_full => outputs_full_140097941532344
        );
        
        core_inst_140097941532400: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941532400,
            fifo_full => fifo_full_140097941532400,
            outputs => outputs_140097941532400,
            outputs_full => outputs_full_140097941532400
        );
        
        core_inst_140097941532456: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941532456,
            fifo_full => fifo_full_140097941532456,
            outputs => outputs_140097941532456,
            outputs_full => outputs_full_140097941532456
        );
        
        core_inst_140097941532512: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941532512,
            fifo_full => fifo_full_140097941532512,
            outputs => outputs_140097941532512,
            outputs_full => outputs_full_140097941532512
        );
        
        core_inst_140097941532568: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941532568,
            fifo_full => fifo_full_140097941532568,
            outputs => outputs_140097941532568,
            outputs_full => outputs_full_140097941532568
        );
        
        core_inst_140097941532624: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941532624,
            fifo_full => fifo_full_140097941532624,
            outputs => outputs_140097941532624,
            outputs_full => outputs_full_140097941532624
        );
        
        core_inst_140097941540936: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941540936,
            fifo_full => fifo_full_140097941540936,
            outputs => outputs_140097941540936,
            outputs_full => outputs_full_140097941540936
        );
        
        core_inst_140097941540992: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941540992,
            fifo_full => fifo_full_140097941540992,
            outputs => outputs_140097941540992,
            outputs_full => outputs_full_140097941540992
        );
        
        core_inst_140097941541048: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941541048,
            fifo_full => fifo_full_140097941541048,
            outputs => outputs_140097941541048,
            outputs_full => outputs_full_140097941541048
        );
        
        core_inst_140097941541104: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941541104,
            fifo_full => fifo_full_140097941541104,
            outputs => outputs_140097941541104,
            outputs_full => outputs_full_140097941541104
        );
        
        core_inst_140097941541160: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941541160,
            fifo_full => fifo_full_140097941541160,
            outputs => outputs_140097941541160,
            outputs_full => outputs_full_140097941541160
        );
        
        core_inst_140097941541216: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941541216,
            fifo_full => fifo_full_140097941541216,
            outputs => outputs_140097941541216,
            outputs_full => outputs_full_140097941541216
        );
        
        core_inst_140097941541272: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941541272,
            fifo_full => fifo_full_140097941541272,
            outputs => outputs_140097941541272,
            outputs_full => outputs_full_140097941541272
        );
        
        core_inst_140097941541328: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941541328,
            fifo_full => fifo_full_140097941541328,
            outputs => outputs_140097941541328,
            outputs_full => outputs_full_140097941541328
        );
        
        core_inst_140097941541384: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941541384,
            fifo_full => fifo_full_140097941541384,
            outputs => outputs_140097941541384,
            outputs_full => outputs_full_140097941541384
        );
        
        core_inst_140097941541440: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941541440,
            fifo_full => fifo_full_140097941541440,
            outputs => outputs_140097941541440,
            outputs_full => outputs_full_140097941541440
        );
        
        core_inst_140097941541496: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941541496,
            fifo_full => fifo_full_140097941541496,
            outputs => outputs_140097941541496,
            outputs_full => outputs_full_140097941541496
        );
        
        core_inst_140097941541552: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941541552,
            fifo_full => fifo_full_140097941541552,
            outputs => outputs_140097941541552,
            outputs_full => outputs_full_140097941541552
        );
        
        core_inst_140097941541608: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941541608,
            fifo_full => fifo_full_140097941541608,
            outputs => outputs_140097941541608,
            outputs_full => outputs_full_140097941541608
        );
        
        core_inst_140097941541664: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941541664,
            fifo_full => fifo_full_140097941541664,
            outputs => outputs_140097941541664,
            outputs_full => outputs_full_140097941541664
        );
        
        core_inst_140097941541720: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941541720,
            fifo_full => fifo_full_140097941541720,
            outputs => outputs_140097941541720,
            outputs_full => outputs_full_140097941541720
        );
        
        core_inst_140097941541776: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941541776,
            fifo_full => fifo_full_140097941541776,
            outputs => outputs_140097941541776,
            outputs_full => outputs_full_140097941541776
        );
        
        core_inst_140097941541832: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941541832,
            fifo_full => fifo_full_140097941541832,
            outputs => outputs_140097941541832,
            outputs_full => outputs_full_140097941541832
        );
        
        core_inst_140097941541888: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941541888,
            fifo_full => fifo_full_140097941541888,
            outputs => outputs_140097941541888,
            outputs_full => outputs_full_140097941541888
        );
        
        core_inst_140097941541944: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941541944,
            fifo_full => fifo_full_140097941541944,
            outputs => outputs_140097941541944,
            outputs_full => outputs_full_140097941541944
        );
        
        core_inst_140097941542000: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941542000,
            fifo_full => fifo_full_140097941542000,
            outputs => outputs_140097941542000,
            outputs_full => outputs_full_140097941542000
        );
        
        core_inst_140097941542056: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941542056,
            fifo_full => fifo_full_140097941542056,
            outputs => outputs_140097941542056,
            outputs_full => outputs_full_140097941542056
        );
        
        core_inst_140097941542112: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941542112,
            fifo_full => fifo_full_140097941542112,
            outputs => outputs_140097941542112,
            outputs_full => outputs_full_140097941542112
        );
        
        core_inst_140097941542168: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941542168,
            fifo_full => fifo_full_140097941542168,
            outputs => outputs_140097941542168,
            outputs_full => outputs_full_140097941542168
        );
        
        core_inst_140097941542224: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941542224,
            fifo_full => fifo_full_140097941542224,
            outputs => outputs_140097941542224,
            outputs_full => outputs_full_140097941542224
        );
        
        core_inst_140097941542280: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941542280,
            fifo_full => fifo_full_140097941542280,
            outputs => outputs_140097941542280,
            outputs_full => outputs_full_140097941542280
        );
        
        core_inst_140097941542336: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941542336,
            fifo_full => fifo_full_140097941542336,
            outputs => outputs_140097941542336,
            outputs_full => outputs_full_140097941542336
        );
        
        core_inst_140097941542392: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941542392,
            fifo_full => fifo_full_140097941542392,
            outputs => outputs_140097941542392,
            outputs_full => outputs_full_140097941542392
        );
        
        core_inst_140097941542448: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941542448,
            fifo_full => fifo_full_140097941542448,
            outputs => outputs_140097941542448,
            outputs_full => outputs_full_140097941542448
        );
        
        core_inst_140097941542504: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941542504,
            fifo_full => fifo_full_140097941542504,
            outputs => outputs_140097941542504,
            outputs_full => outputs_full_140097941542504
        );
        
        core_inst_140097941542560: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941542560,
            fifo_full => fifo_full_140097941542560,
            outputs => outputs_140097941542560,
            outputs_full => outputs_full_140097941542560
        );
        
        core_inst_140097941542616: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941542616,
            fifo_full => fifo_full_140097941542616,
            outputs => outputs_140097941542616,
            outputs_full => outputs_full_140097941542616
        );
        
        core_inst_140097941542672: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941542672,
            fifo_full => fifo_full_140097941542672,
            outputs => outputs_140097941542672,
            outputs_full => outputs_full_140097941542672
        );
        
        core_inst_140097941542728: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941542728,
            fifo_full => fifo_full_140097941542728,
            outputs => outputs_140097941542728,
            outputs_full => outputs_full_140097941542728
        );
        
        core_inst_140097941542784: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941542784,
            fifo_full => fifo_full_140097941542784,
            outputs => outputs_140097941542784,
            outputs_full => outputs_full_140097941542784
        );
        
        core_inst_140097941542840: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941542840,
            fifo_full => fifo_full_140097941542840,
            outputs => outputs_140097941542840,
            outputs_full => outputs_full_140097941542840
        );
        
        core_inst_140097941542896: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941542896,
            fifo_full => fifo_full_140097941542896,
            outputs => outputs_140097941542896,
            outputs_full => outputs_full_140097941542896
        );
        
        core_inst_140097941542952: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941542952,
            fifo_full => fifo_full_140097941542952,
            outputs => outputs_140097941542952,
            outputs_full => outputs_full_140097941542952
        );
        
        core_inst_140097941543008: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941543008,
            fifo_full => fifo_full_140097941543008,
            outputs => outputs_140097941543008,
            outputs_full => outputs_full_140097941543008
        );
        
        core_inst_140097941543064: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941543064,
            fifo_full => fifo_full_140097941543064,
            outputs => outputs_140097941543064,
            outputs_full => outputs_full_140097941543064
        );
        
        core_inst_140097941543120: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941543120,
            fifo_full => fifo_full_140097941543120,
            outputs => outputs_140097941543120,
            outputs_full => outputs_full_140097941543120
        );
        
        core_inst_140097941543176: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941543176,
            fifo_full => fifo_full_140097941543176,
            outputs => outputs_140097941543176,
            outputs_full => outputs_full_140097941543176
        );
        
        core_inst_140097941543232: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941543232,
            fifo_full => fifo_full_140097941543232,
            outputs => outputs_140097941543232,
            outputs_full => outputs_full_140097941543232
        );
        
        core_inst_140097941543288: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941543288,
            fifo_full => fifo_full_140097941543288,
            outputs => outputs_140097941543288,
            outputs_full => outputs_full_140097941543288
        );
        
        core_inst_140097941543344: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941543344,
            fifo_full => fifo_full_140097941543344,
            outputs => outputs_140097941543344,
            outputs_full => outputs_full_140097941543344
        );
        
        core_inst_140097941543400: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941543400,
            fifo_full => fifo_full_140097941543400,
            outputs => outputs_140097941543400,
            outputs_full => outputs_full_140097941543400
        );
        
        core_inst_140097941543456: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941543456,
            fifo_full => fifo_full_140097941543456,
            outputs => outputs_140097941543456,
            outputs_full => outputs_full_140097941543456
        );
        
        core_inst_140097941543512: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941543512,
            fifo_full => fifo_full_140097941543512,
            outputs => outputs_140097941543512,
            outputs_full => outputs_full_140097941543512
        );
        
        core_inst_140097941543568: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941543568,
            fifo_full => fifo_full_140097941543568,
            outputs => outputs_140097941543568,
            outputs_full => outputs_full_140097941543568
        );
        
        core_inst_140097941543624: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941543624,
            fifo_full => fifo_full_140097941543624,
            outputs => outputs_140097941543624,
            outputs_full => outputs_full_140097941543624
        );
        
        core_inst_140097941543680: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941543680,
            fifo_full => fifo_full_140097941543680,
            outputs => outputs_140097941543680,
            outputs_full => outputs_full_140097941543680
        );
        
        core_inst_140097941543736: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941543736,
            fifo_full => fifo_full_140097941543736,
            outputs => outputs_140097941543736,
            outputs_full => outputs_full_140097941543736
        );
        
        core_inst_140097941543792: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941543792,
            fifo_full => fifo_full_140097941543792,
            outputs => outputs_140097941543792,
            outputs_full => outputs_full_140097941543792
        );
        
        core_inst_140097941543848: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941543848,
            fifo_full => fifo_full_140097941543848,
            outputs => outputs_140097941543848,
            outputs_full => outputs_full_140097941543848
        );
        
        core_inst_140097941543904: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941543904,
            fifo_full => fifo_full_140097941543904,
            outputs => outputs_140097941543904,
            outputs_full => outputs_full_140097941543904
        );
        
        core_inst_140097941543960: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941543960,
            fifo_full => fifo_full_140097941543960,
            outputs => outputs_140097941543960,
            outputs_full => outputs_full_140097941543960
        );
        
        core_inst_140097941544016: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941544016,
            fifo_full => fifo_full_140097941544016,
            outputs => outputs_140097941544016,
            outputs_full => outputs_full_140097941544016
        );
        
        core_inst_140097941544072: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941544072,
            fifo_full => fifo_full_140097941544072,
            outputs => outputs_140097941544072,
            outputs_full => outputs_full_140097941544072
        );
        
        core_inst_140097941544128: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941544128,
            fifo_full => fifo_full_140097941544128,
            outputs => outputs_140097941544128,
            outputs_full => outputs_full_140097941544128
        );
        
        core_inst_140097941544184: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941544184,
            fifo_full => fifo_full_140097941544184,
            outputs => outputs_140097941544184,
            outputs_full => outputs_full_140097941544184
        );
        
        core_inst_140097941544240: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941544240,
            fifo_full => fifo_full_140097941544240,
            outputs => outputs_140097941544240,
            outputs_full => outputs_full_140097941544240
        );
        
        core_inst_140097941544296: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941544296,
            fifo_full => fifo_full_140097941544296,
            outputs => outputs_140097941544296,
            outputs_full => outputs_full_140097941544296
        );
        
        core_inst_140097941544352: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941544352,
            fifo_full => fifo_full_140097941544352,
            outputs => outputs_140097941544352,
            outputs_full => outputs_full_140097941544352
        );
        
        core_inst_140097941544408: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941544408,
            fifo_full => fifo_full_140097941544408,
            outputs => outputs_140097941544408,
            outputs_full => outputs_full_140097941544408
        );
        
        core_inst_140097941544464: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941544464,
            fifo_full => fifo_full_140097941544464,
            outputs => outputs_140097941544464,
            outputs_full => outputs_full_140097941544464
        );
        
        core_inst_140097941544520: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941544520,
            fifo_full => fifo_full_140097941544520,
            outputs => outputs_140097941544520,
            outputs_full => outputs_full_140097941544520
        );
        
        core_inst_140097941544576: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941544576,
            fifo_full => fifo_full_140097941544576,
            outputs => outputs_140097941544576,
            outputs_full => outputs_full_140097941544576
        );
        
        core_inst_140097941544632: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941544632,
            fifo_full => fifo_full_140097941544632,
            outputs => outputs_140097941544632,
            outputs_full => outputs_full_140097941544632
        );
        
        core_inst_140097941544688: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941544688,
            fifo_full => fifo_full_140097941544688,
            outputs => outputs_140097941544688,
            outputs_full => outputs_full_140097941544688
        );
        
        core_inst_140097941544744: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941544744,
            fifo_full => fifo_full_140097941544744,
            outputs => outputs_140097941544744,
            outputs_full => outputs_full_140097941544744
        );
        
        core_inst_140097941544800: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941544800,
            fifo_full => fifo_full_140097941544800,
            outputs => outputs_140097941544800,
            outputs_full => outputs_full_140097941544800
        );
        
        core_inst_140097941544856: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941544856,
            fifo_full => fifo_full_140097941544856,
            outputs => outputs_140097941544856,
            outputs_full => outputs_full_140097941544856
        );
        
        core_inst_140097941544912: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941544912,
            fifo_full => fifo_full_140097941544912,
            outputs => outputs_140097941544912,
            outputs_full => outputs_full_140097941544912
        );
        
        core_inst_140097941553224: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941553224,
            fifo_full => fifo_full_140097941553224,
            outputs => outputs_140097941553224,
            outputs_full => outputs_full_140097941553224
        );
        
        core_inst_140097941553280: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941553280,
            fifo_full => fifo_full_140097941553280,
            outputs => outputs_140097941553280,
            outputs_full => outputs_full_140097941553280
        );
        
        core_inst_140097941553336: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941553336,
            fifo_full => fifo_full_140097941553336,
            outputs => outputs_140097941553336,
            outputs_full => outputs_full_140097941553336
        );
        
        core_inst_140097941553392: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941553392,
            fifo_full => fifo_full_140097941553392,
            outputs => outputs_140097941553392,
            outputs_full => outputs_full_140097941553392
        );
        
        core_inst_140097941553448: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941553448,
            fifo_full => fifo_full_140097941553448,
            outputs => outputs_140097941553448,
            outputs_full => outputs_full_140097941553448
        );
        
        core_inst_140097941553504: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941553504,
            fifo_full => fifo_full_140097941553504,
            outputs => outputs_140097941553504,
            outputs_full => outputs_full_140097941553504
        );
        
        core_inst_140097941553560: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941553560,
            fifo_full => fifo_full_140097941553560,
            outputs => outputs_140097941553560,
            outputs_full => outputs_full_140097941553560
        );
        
        core_inst_140097941553616: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941553616,
            fifo_full => fifo_full_140097941553616,
            outputs => outputs_140097941553616,
            outputs_full => outputs_full_140097941553616
        );
        
        core_inst_140097941553672: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941553672,
            fifo_full => fifo_full_140097941553672,
            outputs => outputs_140097941553672,
            outputs_full => outputs_full_140097941553672
        );
        
        core_inst_140097941553728: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941553728,
            fifo_full => fifo_full_140097941553728,
            outputs => outputs_140097941553728,
            outputs_full => outputs_full_140097941553728
        );
        
        core_inst_140097941553784: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941553784,
            fifo_full => fifo_full_140097941553784,
            outputs => outputs_140097941553784,
            outputs_full => outputs_full_140097941553784
        );
        
        core_inst_140097941553840: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941553840,
            fifo_full => fifo_full_140097941553840,
            outputs => outputs_140097941553840,
            outputs_full => outputs_full_140097941553840
        );
        
        core_inst_140097941553896: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941553896,
            fifo_full => fifo_full_140097941553896,
            outputs => outputs_140097941553896,
            outputs_full => outputs_full_140097941553896
        );
        
        core_inst_140097941553952: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941553952,
            fifo_full => fifo_full_140097941553952,
            outputs => outputs_140097941553952,
            outputs_full => outputs_full_140097941553952
        );
        
        core_inst_140097941554008: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941554008,
            fifo_full => fifo_full_140097941554008,
            outputs => outputs_140097941554008,
            outputs_full => outputs_full_140097941554008
        );
        
        core_inst_140097941554064: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941554064,
            fifo_full => fifo_full_140097941554064,
            outputs => outputs_140097941554064,
            outputs_full => outputs_full_140097941554064
        );
        
        core_inst_140097941554120: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941554120,
            fifo_full => fifo_full_140097941554120,
            outputs => outputs_140097941554120,
            outputs_full => outputs_full_140097941554120
        );
        
        core_inst_140097941554176: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941554176,
            fifo_full => fifo_full_140097941554176,
            outputs => outputs_140097941554176,
            outputs_full => outputs_full_140097941554176
        );
        
        core_inst_140097941554232: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941554232,
            fifo_full => fifo_full_140097941554232,
            outputs => outputs_140097941554232,
            outputs_full => outputs_full_140097941554232
        );
        
        core_inst_140097941554288: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941554288,
            fifo_full => fifo_full_140097941554288,
            outputs => outputs_140097941554288,
            outputs_full => outputs_full_140097941554288
        );
        
        core_inst_140097941554344: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941554344,
            fifo_full => fifo_full_140097941554344,
            outputs => outputs_140097941554344,
            outputs_full => outputs_full_140097941554344
        );
        
        core_inst_140097941554400: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941554400,
            fifo_full => fifo_full_140097941554400,
            outputs => outputs_140097941554400,
            outputs_full => outputs_full_140097941554400
        );
        
        core_inst_140097941554456: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941554456,
            fifo_full => fifo_full_140097941554456,
            outputs => outputs_140097941554456,
            outputs_full => outputs_full_140097941554456
        );
        
        core_inst_140097941554512: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941554512,
            fifo_full => fifo_full_140097941554512,
            outputs => outputs_140097941554512,
            outputs_full => outputs_full_140097941554512
        );
        
        core_inst_140097941554568: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941554568,
            fifo_full => fifo_full_140097941554568,
            outputs => outputs_140097941554568,
            outputs_full => outputs_full_140097941554568
        );
        
        core_inst_140097941554624: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941554624,
            fifo_full => fifo_full_140097941554624,
            outputs => outputs_140097941554624,
            outputs_full => outputs_full_140097941554624
        );
        
        core_inst_140097941554680: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941554680,
            fifo_full => fifo_full_140097941554680,
            outputs => outputs_140097941554680,
            outputs_full => outputs_full_140097941554680
        );
        
        core_inst_140097941554736: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941554736,
            fifo_full => fifo_full_140097941554736,
            outputs => outputs_140097941554736,
            outputs_full => outputs_full_140097941554736
        );
        
        core_inst_140097941554792: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941554792,
            fifo_full => fifo_full_140097941554792,
            outputs => outputs_140097941554792,
            outputs_full => outputs_full_140097941554792
        );
        
        core_inst_140097941554848: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941554848,
            fifo_full => fifo_full_140097941554848,
            outputs => outputs_140097941554848,
            outputs_full => outputs_full_140097941554848
        );
        
        core_inst_140097941554904: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941554904,
            fifo_full => fifo_full_140097941554904,
            outputs => outputs_140097941554904,
            outputs_full => outputs_full_140097941554904
        );
        
        core_inst_140097941554960: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941554960,
            fifo_full => fifo_full_140097941554960,
            outputs => outputs_140097941554960,
            outputs_full => outputs_full_140097941554960
        );
        
        core_inst_140097941555016: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941555016,
            fifo_full => fifo_full_140097941555016,
            outputs => outputs_140097941555016,
            outputs_full => outputs_full_140097941555016
        );
        
        core_inst_140097941555072: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941555072,
            fifo_full => fifo_full_140097941555072,
            outputs => outputs_140097941555072,
            outputs_full => outputs_full_140097941555072
        );
        
        core_inst_140097941555128: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941555128,
            fifo_full => fifo_full_140097941555128,
            outputs => outputs_140097941555128,
            outputs_full => outputs_full_140097941555128
        );
        
        core_inst_140097941555184: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941555184,
            fifo_full => fifo_full_140097941555184,
            outputs => outputs_140097941555184,
            outputs_full => outputs_full_140097941555184
        );
        
        core_inst_140097941555240: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941555240,
            fifo_full => fifo_full_140097941555240,
            outputs => outputs_140097941555240,
            outputs_full => outputs_full_140097941555240
        );
        
        core_inst_140097941555296: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941555296,
            fifo_full => fifo_full_140097941555296,
            outputs => outputs_140097941555296,
            outputs_full => outputs_full_140097941555296
        );
        
        core_inst_140097941555352: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941555352,
            fifo_full => fifo_full_140097941555352,
            outputs => outputs_140097941555352,
            outputs_full => outputs_full_140097941555352
        );
        
        core_inst_140097941555408: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941555408,
            fifo_full => fifo_full_140097941555408,
            outputs => outputs_140097941555408,
            outputs_full => outputs_full_140097941555408
        );
        
        core_inst_140097941555464: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941555464,
            fifo_full => fifo_full_140097941555464,
            outputs => outputs_140097941555464,
            outputs_full => outputs_full_140097941555464
        );
        
        core_inst_140097941555520: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941555520,
            fifo_full => fifo_full_140097941555520,
            outputs => outputs_140097941555520,
            outputs_full => outputs_full_140097941555520
        );
        
        core_inst_140097941555576: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941555576,
            fifo_full => fifo_full_140097941555576,
            outputs => outputs_140097941555576,
            outputs_full => outputs_full_140097941555576
        );
        
        core_inst_140097941555632: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941555632,
            fifo_full => fifo_full_140097941555632,
            outputs => outputs_140097941555632,
            outputs_full => outputs_full_140097941555632
        );
        
        core_inst_140097941555688: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140097941555688,
            fifo_full => fifo_full_140097941555688,
            outputs => outputs_140097941555688,
            outputs_full => outputs_full_140097941555688
        );
        
        outputs <= outputs_140097941555688;
        outputs_full_140097941555688 <= outputs_full;

end behav;

