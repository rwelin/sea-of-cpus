
library ieee;
use ieee.std_logic_1164.all;
use work.core_config.all;
use work.all;

entity Grid8 is
    port (
        clk: in std_logic;
        clk_en: in std_logic;
        reset: in std_logic;
        addr: in ram_addr;
        data: in word;
        we: in std_logic;
        fifo_inputs: in core_fifo_inputs_t;
        fifo_full: out std_logic_vector(0 to NUM_CORE_FIFOS-1);
        outputs: out core_fifo_inputs_t;
        outputs_full: in std_logic_vector(0 to NUM_CORE_FIFOS-1)
    );
end Grid8;

architecture behav of Grid8 is

    
        signal fifo_inputs_140108714687736: core_fifo_inputs_t;
        signal fifo_full_140108714687736: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714687736: core_fifo_inputs_t;
        signal outputs_full_140108714687736: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714687960: core_fifo_inputs_t;
        signal fifo_full_140108714687960: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714687960: core_fifo_inputs_t;
        signal outputs_full_140108714687960: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714687904: core_fifo_inputs_t;
        signal fifo_full_140108714687904: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714687904: core_fifo_inputs_t;
        signal outputs_full_140108714687904: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714688016: core_fifo_inputs_t;
        signal fifo_full_140108714688016: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714688016: core_fifo_inputs_t;
        signal outputs_full_140108714688016: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714688072: core_fifo_inputs_t;
        signal fifo_full_140108714688072: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714688072: core_fifo_inputs_t;
        signal outputs_full_140108714688072: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714688128: core_fifo_inputs_t;
        signal fifo_full_140108714688128: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714688128: core_fifo_inputs_t;
        signal outputs_full_140108714688128: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714688184: core_fifo_inputs_t;
        signal fifo_full_140108714688184: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714688184: core_fifo_inputs_t;
        signal outputs_full_140108714688184: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714688240: core_fifo_inputs_t;
        signal fifo_full_140108714688240: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714688240: core_fifo_inputs_t;
        signal outputs_full_140108714688240: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714688296: core_fifo_inputs_t;
        signal fifo_full_140108714688296: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714688296: core_fifo_inputs_t;
        signal outputs_full_140108714688296: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714687848: core_fifo_inputs_t;
        signal fifo_full_140108714687848: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714687848: core_fifo_inputs_t;
        signal outputs_full_140108714687848: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714688352: core_fifo_inputs_t;
        signal fifo_full_140108714688352: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714688352: core_fifo_inputs_t;
        signal outputs_full_140108714688352: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714688408: core_fifo_inputs_t;
        signal fifo_full_140108714688408: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714688408: core_fifo_inputs_t;
        signal outputs_full_140108714688408: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714688464: core_fifo_inputs_t;
        signal fifo_full_140108714688464: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714688464: core_fifo_inputs_t;
        signal outputs_full_140108714688464: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714733640: core_fifo_inputs_t;
        signal fifo_full_140108714733640: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714733640: core_fifo_inputs_t;
        signal outputs_full_140108714733640: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714733696: core_fifo_inputs_t;
        signal fifo_full_140108714733696: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714733696: core_fifo_inputs_t;
        signal outputs_full_140108714733696: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714733752: core_fifo_inputs_t;
        signal fifo_full_140108714733752: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714733752: core_fifo_inputs_t;
        signal outputs_full_140108714733752: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714733808: core_fifo_inputs_t;
        signal fifo_full_140108714733808: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714733808: core_fifo_inputs_t;
        signal outputs_full_140108714733808: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714733864: core_fifo_inputs_t;
        signal fifo_full_140108714733864: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714733864: core_fifo_inputs_t;
        signal outputs_full_140108714733864: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714733920: core_fifo_inputs_t;
        signal fifo_full_140108714733920: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714733920: core_fifo_inputs_t;
        signal outputs_full_140108714733920: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714733976: core_fifo_inputs_t;
        signal fifo_full_140108714733976: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714733976: core_fifo_inputs_t;
        signal outputs_full_140108714733976: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714734032: core_fifo_inputs_t;
        signal fifo_full_140108714734032: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714734032: core_fifo_inputs_t;
        signal outputs_full_140108714734032: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714734088: core_fifo_inputs_t;
        signal fifo_full_140108714734088: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714734088: core_fifo_inputs_t;
        signal outputs_full_140108714734088: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714734144: core_fifo_inputs_t;
        signal fifo_full_140108714734144: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714734144: core_fifo_inputs_t;
        signal outputs_full_140108714734144: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714734200: core_fifo_inputs_t;
        signal fifo_full_140108714734200: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714734200: core_fifo_inputs_t;
        signal outputs_full_140108714734200: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714734256: core_fifo_inputs_t;
        signal fifo_full_140108714734256: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714734256: core_fifo_inputs_t;
        signal outputs_full_140108714734256: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714734312: core_fifo_inputs_t;
        signal fifo_full_140108714734312: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714734312: core_fifo_inputs_t;
        signal outputs_full_140108714734312: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714734368: core_fifo_inputs_t;
        signal fifo_full_140108714734368: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714734368: core_fifo_inputs_t;
        signal outputs_full_140108714734368: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714734424: core_fifo_inputs_t;
        signal fifo_full_140108714734424: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714734424: core_fifo_inputs_t;
        signal outputs_full_140108714734424: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714734480: core_fifo_inputs_t;
        signal fifo_full_140108714734480: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714734480: core_fifo_inputs_t;
        signal outputs_full_140108714734480: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714734536: core_fifo_inputs_t;
        signal fifo_full_140108714734536: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714734536: core_fifo_inputs_t;
        signal outputs_full_140108714734536: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714734592: core_fifo_inputs_t;
        signal fifo_full_140108714734592: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714734592: core_fifo_inputs_t;
        signal outputs_full_140108714734592: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714734648: core_fifo_inputs_t;
        signal fifo_full_140108714734648: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714734648: core_fifo_inputs_t;
        signal outputs_full_140108714734648: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714734704: core_fifo_inputs_t;
        signal fifo_full_140108714734704: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714734704: core_fifo_inputs_t;
        signal outputs_full_140108714734704: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714734760: core_fifo_inputs_t;
        signal fifo_full_140108714734760: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714734760: core_fifo_inputs_t;
        signal outputs_full_140108714734760: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714734816: core_fifo_inputs_t;
        signal fifo_full_140108714734816: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714734816: core_fifo_inputs_t;
        signal outputs_full_140108714734816: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714734872: core_fifo_inputs_t;
        signal fifo_full_140108714734872: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714734872: core_fifo_inputs_t;
        signal outputs_full_140108714734872: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714734928: core_fifo_inputs_t;
        signal fifo_full_140108714734928: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714734928: core_fifo_inputs_t;
        signal outputs_full_140108714734928: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714734984: core_fifo_inputs_t;
        signal fifo_full_140108714734984: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714734984: core_fifo_inputs_t;
        signal outputs_full_140108714734984: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714735040: core_fifo_inputs_t;
        signal fifo_full_140108714735040: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714735040: core_fifo_inputs_t;
        signal outputs_full_140108714735040: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714735096: core_fifo_inputs_t;
        signal fifo_full_140108714735096: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714735096: core_fifo_inputs_t;
        signal outputs_full_140108714735096: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714735152: core_fifo_inputs_t;
        signal fifo_full_140108714735152: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714735152: core_fifo_inputs_t;
        signal outputs_full_140108714735152: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714735208: core_fifo_inputs_t;
        signal fifo_full_140108714735208: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714735208: core_fifo_inputs_t;
        signal outputs_full_140108714735208: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714735264: core_fifo_inputs_t;
        signal fifo_full_140108714735264: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714735264: core_fifo_inputs_t;
        signal outputs_full_140108714735264: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714735320: core_fifo_inputs_t;
        signal fifo_full_140108714735320: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714735320: core_fifo_inputs_t;
        signal outputs_full_140108714735320: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714735376: core_fifo_inputs_t;
        signal fifo_full_140108714735376: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714735376: core_fifo_inputs_t;
        signal outputs_full_140108714735376: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714735432: core_fifo_inputs_t;
        signal fifo_full_140108714735432: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714735432: core_fifo_inputs_t;
        signal outputs_full_140108714735432: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714735488: core_fifo_inputs_t;
        signal fifo_full_140108714735488: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714735488: core_fifo_inputs_t;
        signal outputs_full_140108714735488: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714735544: core_fifo_inputs_t;
        signal fifo_full_140108714735544: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714735544: core_fifo_inputs_t;
        signal outputs_full_140108714735544: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714735600: core_fifo_inputs_t;
        signal fifo_full_140108714735600: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714735600: core_fifo_inputs_t;
        signal outputs_full_140108714735600: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714735656: core_fifo_inputs_t;
        signal fifo_full_140108714735656: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714735656: core_fifo_inputs_t;
        signal outputs_full_140108714735656: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714735712: core_fifo_inputs_t;
        signal fifo_full_140108714735712: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714735712: core_fifo_inputs_t;
        signal outputs_full_140108714735712: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714735768: core_fifo_inputs_t;
        signal fifo_full_140108714735768: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714735768: core_fifo_inputs_t;
        signal outputs_full_140108714735768: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714735824: core_fifo_inputs_t;
        signal fifo_full_140108714735824: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714735824: core_fifo_inputs_t;
        signal outputs_full_140108714735824: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714735880: core_fifo_inputs_t;
        signal fifo_full_140108714735880: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714735880: core_fifo_inputs_t;
        signal outputs_full_140108714735880: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714735936: core_fifo_inputs_t;
        signal fifo_full_140108714735936: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714735936: core_fifo_inputs_t;
        signal outputs_full_140108714735936: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714735992: core_fifo_inputs_t;
        signal fifo_full_140108714735992: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714735992: core_fifo_inputs_t;
        signal outputs_full_140108714735992: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714736048: core_fifo_inputs_t;
        signal fifo_full_140108714736048: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714736048: core_fifo_inputs_t;
        signal outputs_full_140108714736048: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714736104: core_fifo_inputs_t;
        signal fifo_full_140108714736104: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714736104: core_fifo_inputs_t;
        signal outputs_full_140108714736104: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714736160: core_fifo_inputs_t;
        signal fifo_full_140108714736160: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714736160: core_fifo_inputs_t;
        signal outputs_full_140108714736160: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714736216: core_fifo_inputs_t;
        signal fifo_full_140108714736216: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714736216: core_fifo_inputs_t;
        signal outputs_full_140108714736216: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714736272: core_fifo_inputs_t;
        signal fifo_full_140108714736272: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714736272: core_fifo_inputs_t;
        signal outputs_full_140108714736272: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714736328: core_fifo_inputs_t;
        signal fifo_full_140108714736328: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714736328: core_fifo_inputs_t;
        signal outputs_full_140108714736328: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714736384: core_fifo_inputs_t;
        signal fifo_full_140108714736384: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714736384: core_fifo_inputs_t;
        signal outputs_full_140108714736384: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140108714736440: core_fifo_inputs_t;
        signal fifo_full_140108714736440: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140108714736440: core_fifo_inputs_t;
        signal outputs_full_140108714736440: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        

begin

        outputs(0) <= outputs_140108714736440(0);
        outputs_full_140108714736440(0) <= outputs_full(0);

        fifo_inputs_140108714687736(1) <= fifo_inputs(1);
        fifo_full(1) <= fifo_full_140108714687736(1);
    
        fifo_inputs_140108714687960(1) <= outputs_140108714687736(0);
        outputs_full_140108714687736(0) <= fifo_full_140108714687960(1);
        
        fifo_inputs_140108714688296(3) <= outputs_140108714687736(2);
        outputs_full_140108714687736(2) <= fifo_full_140108714688296(3);
        
        fifo_inputs_140108714687904(1) <= outputs_140108714687960(0);
        outputs_full_140108714687960(0) <= fifo_full_140108714687904(1);
        
        fifo_inputs_140108714687736(0) <= outputs_140108714687960(1);
        outputs_full_140108714687960(1) <= fifo_full_140108714687736(0);
        
        fifo_inputs_140108714687848(3) <= outputs_140108714687960(2);
        outputs_full_140108714687960(2) <= fifo_full_140108714687848(3);
        
        fifo_inputs_140108714688016(1) <= outputs_140108714687904(0);
        outputs_full_140108714687904(0) <= fifo_full_140108714688016(1);
        
        fifo_inputs_140108714687960(0) <= outputs_140108714687904(1);
        outputs_full_140108714687904(1) <= fifo_full_140108714687960(0);
        
        fifo_inputs_140108714688352(3) <= outputs_140108714687904(2);
        outputs_full_140108714687904(2) <= fifo_full_140108714688352(3);
        
        fifo_inputs_140108714688072(1) <= outputs_140108714688016(0);
        outputs_full_140108714688016(0) <= fifo_full_140108714688072(1);
        
        fifo_inputs_140108714687904(0) <= outputs_140108714688016(1);
        outputs_full_140108714688016(1) <= fifo_full_140108714687904(0);
        
        fifo_inputs_140108714688408(3) <= outputs_140108714688016(2);
        outputs_full_140108714688016(2) <= fifo_full_140108714688408(3);
        
        fifo_inputs_140108714688128(1) <= outputs_140108714688072(0);
        outputs_full_140108714688072(0) <= fifo_full_140108714688128(1);
        
        fifo_inputs_140108714688016(0) <= outputs_140108714688072(1);
        outputs_full_140108714688072(1) <= fifo_full_140108714688016(0);
        
        fifo_inputs_140108714688464(3) <= outputs_140108714688072(2);
        outputs_full_140108714688072(2) <= fifo_full_140108714688464(3);
        
        fifo_inputs_140108714688184(1) <= outputs_140108714688128(0);
        outputs_full_140108714688128(0) <= fifo_full_140108714688184(1);
        
        fifo_inputs_140108714688072(0) <= outputs_140108714688128(1);
        outputs_full_140108714688128(1) <= fifo_full_140108714688072(0);
        
        fifo_inputs_140108714733640(3) <= outputs_140108714688128(2);
        outputs_full_140108714688128(2) <= fifo_full_140108714733640(3);
        
        fifo_inputs_140108714688240(1) <= outputs_140108714688184(0);
        outputs_full_140108714688184(0) <= fifo_full_140108714688240(1);
        
        fifo_inputs_140108714688128(0) <= outputs_140108714688184(1);
        outputs_full_140108714688184(1) <= fifo_full_140108714688128(0);
        
        fifo_inputs_140108714733696(3) <= outputs_140108714688184(2);
        outputs_full_140108714688184(2) <= fifo_full_140108714733696(3);
        
        fifo_inputs_140108714688184(0) <= outputs_140108714688240(1);
        outputs_full_140108714688240(1) <= fifo_full_140108714688184(0);
        
        fifo_inputs_140108714733752(3) <= outputs_140108714688240(2);
        outputs_full_140108714688240(2) <= fifo_full_140108714733752(3);
        
        fifo_inputs_140108714687848(1) <= outputs_140108714688296(0);
        outputs_full_140108714688296(0) <= fifo_full_140108714687848(1);
        
        fifo_inputs_140108714733808(3) <= outputs_140108714688296(2);
        outputs_full_140108714688296(2) <= fifo_full_140108714733808(3);
        
        fifo_inputs_140108714687736(2) <= outputs_140108714688296(3);
        outputs_full_140108714688296(3) <= fifo_full_140108714687736(2);
        
        fifo_inputs_140108714688352(1) <= outputs_140108714687848(0);
        outputs_full_140108714687848(0) <= fifo_full_140108714688352(1);
        
        fifo_inputs_140108714688296(0) <= outputs_140108714687848(1);
        outputs_full_140108714687848(1) <= fifo_full_140108714688296(0);
        
        fifo_inputs_140108714733864(3) <= outputs_140108714687848(2);
        outputs_full_140108714687848(2) <= fifo_full_140108714733864(3);
        
        fifo_inputs_140108714687960(2) <= outputs_140108714687848(3);
        outputs_full_140108714687848(3) <= fifo_full_140108714687960(2);
        
        fifo_inputs_140108714688408(1) <= outputs_140108714688352(0);
        outputs_full_140108714688352(0) <= fifo_full_140108714688408(1);
        
        fifo_inputs_140108714687848(0) <= outputs_140108714688352(1);
        outputs_full_140108714688352(1) <= fifo_full_140108714687848(0);
        
        fifo_inputs_140108714733920(3) <= outputs_140108714688352(2);
        outputs_full_140108714688352(2) <= fifo_full_140108714733920(3);
        
        fifo_inputs_140108714687904(2) <= outputs_140108714688352(3);
        outputs_full_140108714688352(3) <= fifo_full_140108714687904(2);
        
        fifo_inputs_140108714688464(1) <= outputs_140108714688408(0);
        outputs_full_140108714688408(0) <= fifo_full_140108714688464(1);
        
        fifo_inputs_140108714688352(0) <= outputs_140108714688408(1);
        outputs_full_140108714688408(1) <= fifo_full_140108714688352(0);
        
        fifo_inputs_140108714733976(3) <= outputs_140108714688408(2);
        outputs_full_140108714688408(2) <= fifo_full_140108714733976(3);
        
        fifo_inputs_140108714688016(2) <= outputs_140108714688408(3);
        outputs_full_140108714688408(3) <= fifo_full_140108714688016(2);
        
        fifo_inputs_140108714733640(1) <= outputs_140108714688464(0);
        outputs_full_140108714688464(0) <= fifo_full_140108714733640(1);
        
        fifo_inputs_140108714688408(0) <= outputs_140108714688464(1);
        outputs_full_140108714688464(1) <= fifo_full_140108714688408(0);
        
        fifo_inputs_140108714734032(3) <= outputs_140108714688464(2);
        outputs_full_140108714688464(2) <= fifo_full_140108714734032(3);
        
        fifo_inputs_140108714688072(2) <= outputs_140108714688464(3);
        outputs_full_140108714688464(3) <= fifo_full_140108714688072(2);
        
        fifo_inputs_140108714733696(1) <= outputs_140108714733640(0);
        outputs_full_140108714733640(0) <= fifo_full_140108714733696(1);
        
        fifo_inputs_140108714688464(0) <= outputs_140108714733640(1);
        outputs_full_140108714733640(1) <= fifo_full_140108714688464(0);
        
        fifo_inputs_140108714734088(3) <= outputs_140108714733640(2);
        outputs_full_140108714733640(2) <= fifo_full_140108714734088(3);
        
        fifo_inputs_140108714688128(2) <= outputs_140108714733640(3);
        outputs_full_140108714733640(3) <= fifo_full_140108714688128(2);
        
        fifo_inputs_140108714733752(1) <= outputs_140108714733696(0);
        outputs_full_140108714733696(0) <= fifo_full_140108714733752(1);
        
        fifo_inputs_140108714733640(0) <= outputs_140108714733696(1);
        outputs_full_140108714733696(1) <= fifo_full_140108714733640(0);
        
        fifo_inputs_140108714734144(3) <= outputs_140108714733696(2);
        outputs_full_140108714733696(2) <= fifo_full_140108714734144(3);
        
        fifo_inputs_140108714688184(2) <= outputs_140108714733696(3);
        outputs_full_140108714733696(3) <= fifo_full_140108714688184(2);
        
        fifo_inputs_140108714733696(0) <= outputs_140108714733752(1);
        outputs_full_140108714733752(1) <= fifo_full_140108714733696(0);
        
        fifo_inputs_140108714734200(3) <= outputs_140108714733752(2);
        outputs_full_140108714733752(2) <= fifo_full_140108714734200(3);
        
        fifo_inputs_140108714688240(2) <= outputs_140108714733752(3);
        outputs_full_140108714733752(3) <= fifo_full_140108714688240(2);
        
        fifo_inputs_140108714733864(1) <= outputs_140108714733808(0);
        outputs_full_140108714733808(0) <= fifo_full_140108714733864(1);
        
        fifo_inputs_140108714734256(3) <= outputs_140108714733808(2);
        outputs_full_140108714733808(2) <= fifo_full_140108714734256(3);
        
        fifo_inputs_140108714688296(2) <= outputs_140108714733808(3);
        outputs_full_140108714733808(3) <= fifo_full_140108714688296(2);
        
        fifo_inputs_140108714733920(1) <= outputs_140108714733864(0);
        outputs_full_140108714733864(0) <= fifo_full_140108714733920(1);
        
        fifo_inputs_140108714733808(0) <= outputs_140108714733864(1);
        outputs_full_140108714733864(1) <= fifo_full_140108714733808(0);
        
        fifo_inputs_140108714734312(3) <= outputs_140108714733864(2);
        outputs_full_140108714733864(2) <= fifo_full_140108714734312(3);
        
        fifo_inputs_140108714687848(2) <= outputs_140108714733864(3);
        outputs_full_140108714733864(3) <= fifo_full_140108714687848(2);
        
        fifo_inputs_140108714733976(1) <= outputs_140108714733920(0);
        outputs_full_140108714733920(0) <= fifo_full_140108714733976(1);
        
        fifo_inputs_140108714733864(0) <= outputs_140108714733920(1);
        outputs_full_140108714733920(1) <= fifo_full_140108714733864(0);
        
        fifo_inputs_140108714734368(3) <= outputs_140108714733920(2);
        outputs_full_140108714733920(2) <= fifo_full_140108714734368(3);
        
        fifo_inputs_140108714688352(2) <= outputs_140108714733920(3);
        outputs_full_140108714733920(3) <= fifo_full_140108714688352(2);
        
        fifo_inputs_140108714734032(1) <= outputs_140108714733976(0);
        outputs_full_140108714733976(0) <= fifo_full_140108714734032(1);
        
        fifo_inputs_140108714733920(0) <= outputs_140108714733976(1);
        outputs_full_140108714733976(1) <= fifo_full_140108714733920(0);
        
        fifo_inputs_140108714734424(3) <= outputs_140108714733976(2);
        outputs_full_140108714733976(2) <= fifo_full_140108714734424(3);
        
        fifo_inputs_140108714688408(2) <= outputs_140108714733976(3);
        outputs_full_140108714733976(3) <= fifo_full_140108714688408(2);
        
        fifo_inputs_140108714734088(1) <= outputs_140108714734032(0);
        outputs_full_140108714734032(0) <= fifo_full_140108714734088(1);
        
        fifo_inputs_140108714733976(0) <= outputs_140108714734032(1);
        outputs_full_140108714734032(1) <= fifo_full_140108714733976(0);
        
        fifo_inputs_140108714734480(3) <= outputs_140108714734032(2);
        outputs_full_140108714734032(2) <= fifo_full_140108714734480(3);
        
        fifo_inputs_140108714688464(2) <= outputs_140108714734032(3);
        outputs_full_140108714734032(3) <= fifo_full_140108714688464(2);
        
        fifo_inputs_140108714734144(1) <= outputs_140108714734088(0);
        outputs_full_140108714734088(0) <= fifo_full_140108714734144(1);
        
        fifo_inputs_140108714734032(0) <= outputs_140108714734088(1);
        outputs_full_140108714734088(1) <= fifo_full_140108714734032(0);
        
        fifo_inputs_140108714734536(3) <= outputs_140108714734088(2);
        outputs_full_140108714734088(2) <= fifo_full_140108714734536(3);
        
        fifo_inputs_140108714733640(2) <= outputs_140108714734088(3);
        outputs_full_140108714734088(3) <= fifo_full_140108714733640(2);
        
        fifo_inputs_140108714734200(1) <= outputs_140108714734144(0);
        outputs_full_140108714734144(0) <= fifo_full_140108714734200(1);
        
        fifo_inputs_140108714734088(0) <= outputs_140108714734144(1);
        outputs_full_140108714734144(1) <= fifo_full_140108714734088(0);
        
        fifo_inputs_140108714734592(3) <= outputs_140108714734144(2);
        outputs_full_140108714734144(2) <= fifo_full_140108714734592(3);
        
        fifo_inputs_140108714733696(2) <= outputs_140108714734144(3);
        outputs_full_140108714734144(3) <= fifo_full_140108714733696(2);
        
        fifo_inputs_140108714734144(0) <= outputs_140108714734200(1);
        outputs_full_140108714734200(1) <= fifo_full_140108714734144(0);
        
        fifo_inputs_140108714734648(3) <= outputs_140108714734200(2);
        outputs_full_140108714734200(2) <= fifo_full_140108714734648(3);
        
        fifo_inputs_140108714733752(2) <= outputs_140108714734200(3);
        outputs_full_140108714734200(3) <= fifo_full_140108714733752(2);
        
        fifo_inputs_140108714734312(1) <= outputs_140108714734256(0);
        outputs_full_140108714734256(0) <= fifo_full_140108714734312(1);
        
        fifo_inputs_140108714734704(3) <= outputs_140108714734256(2);
        outputs_full_140108714734256(2) <= fifo_full_140108714734704(3);
        
        fifo_inputs_140108714733808(2) <= outputs_140108714734256(3);
        outputs_full_140108714734256(3) <= fifo_full_140108714733808(2);
        
        fifo_inputs_140108714734368(1) <= outputs_140108714734312(0);
        outputs_full_140108714734312(0) <= fifo_full_140108714734368(1);
        
        fifo_inputs_140108714734256(0) <= outputs_140108714734312(1);
        outputs_full_140108714734312(1) <= fifo_full_140108714734256(0);
        
        fifo_inputs_140108714734760(3) <= outputs_140108714734312(2);
        outputs_full_140108714734312(2) <= fifo_full_140108714734760(3);
        
        fifo_inputs_140108714733864(2) <= outputs_140108714734312(3);
        outputs_full_140108714734312(3) <= fifo_full_140108714733864(2);
        
        fifo_inputs_140108714734424(1) <= outputs_140108714734368(0);
        outputs_full_140108714734368(0) <= fifo_full_140108714734424(1);
        
        fifo_inputs_140108714734312(0) <= outputs_140108714734368(1);
        outputs_full_140108714734368(1) <= fifo_full_140108714734312(0);
        
        fifo_inputs_140108714734816(3) <= outputs_140108714734368(2);
        outputs_full_140108714734368(2) <= fifo_full_140108714734816(3);
        
        fifo_inputs_140108714733920(2) <= outputs_140108714734368(3);
        outputs_full_140108714734368(3) <= fifo_full_140108714733920(2);
        
        fifo_inputs_140108714734480(1) <= outputs_140108714734424(0);
        outputs_full_140108714734424(0) <= fifo_full_140108714734480(1);
        
        fifo_inputs_140108714734368(0) <= outputs_140108714734424(1);
        outputs_full_140108714734424(1) <= fifo_full_140108714734368(0);
        
        fifo_inputs_140108714734872(3) <= outputs_140108714734424(2);
        outputs_full_140108714734424(2) <= fifo_full_140108714734872(3);
        
        fifo_inputs_140108714733976(2) <= outputs_140108714734424(3);
        outputs_full_140108714734424(3) <= fifo_full_140108714733976(2);
        
        fifo_inputs_140108714734536(1) <= outputs_140108714734480(0);
        outputs_full_140108714734480(0) <= fifo_full_140108714734536(1);
        
        fifo_inputs_140108714734424(0) <= outputs_140108714734480(1);
        outputs_full_140108714734480(1) <= fifo_full_140108714734424(0);
        
        fifo_inputs_140108714734928(3) <= outputs_140108714734480(2);
        outputs_full_140108714734480(2) <= fifo_full_140108714734928(3);
        
        fifo_inputs_140108714734032(2) <= outputs_140108714734480(3);
        outputs_full_140108714734480(3) <= fifo_full_140108714734032(2);
        
        fifo_inputs_140108714734592(1) <= outputs_140108714734536(0);
        outputs_full_140108714734536(0) <= fifo_full_140108714734592(1);
        
        fifo_inputs_140108714734480(0) <= outputs_140108714734536(1);
        outputs_full_140108714734536(1) <= fifo_full_140108714734480(0);
        
        fifo_inputs_140108714734984(3) <= outputs_140108714734536(2);
        outputs_full_140108714734536(2) <= fifo_full_140108714734984(3);
        
        fifo_inputs_140108714734088(2) <= outputs_140108714734536(3);
        outputs_full_140108714734536(3) <= fifo_full_140108714734088(2);
        
        fifo_inputs_140108714734648(1) <= outputs_140108714734592(0);
        outputs_full_140108714734592(0) <= fifo_full_140108714734648(1);
        
        fifo_inputs_140108714734536(0) <= outputs_140108714734592(1);
        outputs_full_140108714734592(1) <= fifo_full_140108714734536(0);
        
        fifo_inputs_140108714735040(3) <= outputs_140108714734592(2);
        outputs_full_140108714734592(2) <= fifo_full_140108714735040(3);
        
        fifo_inputs_140108714734144(2) <= outputs_140108714734592(3);
        outputs_full_140108714734592(3) <= fifo_full_140108714734144(2);
        
        fifo_inputs_140108714734592(0) <= outputs_140108714734648(1);
        outputs_full_140108714734648(1) <= fifo_full_140108714734592(0);
        
        fifo_inputs_140108714735096(3) <= outputs_140108714734648(2);
        outputs_full_140108714734648(2) <= fifo_full_140108714735096(3);
        
        fifo_inputs_140108714734200(2) <= outputs_140108714734648(3);
        outputs_full_140108714734648(3) <= fifo_full_140108714734200(2);
        
        fifo_inputs_140108714734760(1) <= outputs_140108714734704(0);
        outputs_full_140108714734704(0) <= fifo_full_140108714734760(1);
        
        fifo_inputs_140108714735152(3) <= outputs_140108714734704(2);
        outputs_full_140108714734704(2) <= fifo_full_140108714735152(3);
        
        fifo_inputs_140108714734256(2) <= outputs_140108714734704(3);
        outputs_full_140108714734704(3) <= fifo_full_140108714734256(2);
        
        fifo_inputs_140108714734816(1) <= outputs_140108714734760(0);
        outputs_full_140108714734760(0) <= fifo_full_140108714734816(1);
        
        fifo_inputs_140108714734704(0) <= outputs_140108714734760(1);
        outputs_full_140108714734760(1) <= fifo_full_140108714734704(0);
        
        fifo_inputs_140108714735208(3) <= outputs_140108714734760(2);
        outputs_full_140108714734760(2) <= fifo_full_140108714735208(3);
        
        fifo_inputs_140108714734312(2) <= outputs_140108714734760(3);
        outputs_full_140108714734760(3) <= fifo_full_140108714734312(2);
        
        fifo_inputs_140108714734872(1) <= outputs_140108714734816(0);
        outputs_full_140108714734816(0) <= fifo_full_140108714734872(1);
        
        fifo_inputs_140108714734760(0) <= outputs_140108714734816(1);
        outputs_full_140108714734816(1) <= fifo_full_140108714734760(0);
        
        fifo_inputs_140108714735264(3) <= outputs_140108714734816(2);
        outputs_full_140108714734816(2) <= fifo_full_140108714735264(3);
        
        fifo_inputs_140108714734368(2) <= outputs_140108714734816(3);
        outputs_full_140108714734816(3) <= fifo_full_140108714734368(2);
        
        fifo_inputs_140108714734928(1) <= outputs_140108714734872(0);
        outputs_full_140108714734872(0) <= fifo_full_140108714734928(1);
        
        fifo_inputs_140108714734816(0) <= outputs_140108714734872(1);
        outputs_full_140108714734872(1) <= fifo_full_140108714734816(0);
        
        fifo_inputs_140108714735320(3) <= outputs_140108714734872(2);
        outputs_full_140108714734872(2) <= fifo_full_140108714735320(3);
        
        fifo_inputs_140108714734424(2) <= outputs_140108714734872(3);
        outputs_full_140108714734872(3) <= fifo_full_140108714734424(2);
        
        fifo_inputs_140108714734984(1) <= outputs_140108714734928(0);
        outputs_full_140108714734928(0) <= fifo_full_140108714734984(1);
        
        fifo_inputs_140108714734872(0) <= outputs_140108714734928(1);
        outputs_full_140108714734928(1) <= fifo_full_140108714734872(0);
        
        fifo_inputs_140108714735376(3) <= outputs_140108714734928(2);
        outputs_full_140108714734928(2) <= fifo_full_140108714735376(3);
        
        fifo_inputs_140108714734480(2) <= outputs_140108714734928(3);
        outputs_full_140108714734928(3) <= fifo_full_140108714734480(2);
        
        fifo_inputs_140108714735040(1) <= outputs_140108714734984(0);
        outputs_full_140108714734984(0) <= fifo_full_140108714735040(1);
        
        fifo_inputs_140108714734928(0) <= outputs_140108714734984(1);
        outputs_full_140108714734984(1) <= fifo_full_140108714734928(0);
        
        fifo_inputs_140108714735432(3) <= outputs_140108714734984(2);
        outputs_full_140108714734984(2) <= fifo_full_140108714735432(3);
        
        fifo_inputs_140108714734536(2) <= outputs_140108714734984(3);
        outputs_full_140108714734984(3) <= fifo_full_140108714734536(2);
        
        fifo_inputs_140108714735096(1) <= outputs_140108714735040(0);
        outputs_full_140108714735040(0) <= fifo_full_140108714735096(1);
        
        fifo_inputs_140108714734984(0) <= outputs_140108714735040(1);
        outputs_full_140108714735040(1) <= fifo_full_140108714734984(0);
        
        fifo_inputs_140108714735488(3) <= outputs_140108714735040(2);
        outputs_full_140108714735040(2) <= fifo_full_140108714735488(3);
        
        fifo_inputs_140108714734592(2) <= outputs_140108714735040(3);
        outputs_full_140108714735040(3) <= fifo_full_140108714734592(2);
        
        fifo_inputs_140108714735040(0) <= outputs_140108714735096(1);
        outputs_full_140108714735096(1) <= fifo_full_140108714735040(0);
        
        fifo_inputs_140108714735544(3) <= outputs_140108714735096(2);
        outputs_full_140108714735096(2) <= fifo_full_140108714735544(3);
        
        fifo_inputs_140108714734648(2) <= outputs_140108714735096(3);
        outputs_full_140108714735096(3) <= fifo_full_140108714734648(2);
        
        fifo_inputs_140108714735208(1) <= outputs_140108714735152(0);
        outputs_full_140108714735152(0) <= fifo_full_140108714735208(1);
        
        fifo_inputs_140108714735600(3) <= outputs_140108714735152(2);
        outputs_full_140108714735152(2) <= fifo_full_140108714735600(3);
        
        fifo_inputs_140108714734704(2) <= outputs_140108714735152(3);
        outputs_full_140108714735152(3) <= fifo_full_140108714734704(2);
        
        fifo_inputs_140108714735264(1) <= outputs_140108714735208(0);
        outputs_full_140108714735208(0) <= fifo_full_140108714735264(1);
        
        fifo_inputs_140108714735152(0) <= outputs_140108714735208(1);
        outputs_full_140108714735208(1) <= fifo_full_140108714735152(0);
        
        fifo_inputs_140108714735656(3) <= outputs_140108714735208(2);
        outputs_full_140108714735208(2) <= fifo_full_140108714735656(3);
        
        fifo_inputs_140108714734760(2) <= outputs_140108714735208(3);
        outputs_full_140108714735208(3) <= fifo_full_140108714734760(2);
        
        fifo_inputs_140108714735320(1) <= outputs_140108714735264(0);
        outputs_full_140108714735264(0) <= fifo_full_140108714735320(1);
        
        fifo_inputs_140108714735208(0) <= outputs_140108714735264(1);
        outputs_full_140108714735264(1) <= fifo_full_140108714735208(0);
        
        fifo_inputs_140108714735712(3) <= outputs_140108714735264(2);
        outputs_full_140108714735264(2) <= fifo_full_140108714735712(3);
        
        fifo_inputs_140108714734816(2) <= outputs_140108714735264(3);
        outputs_full_140108714735264(3) <= fifo_full_140108714734816(2);
        
        fifo_inputs_140108714735376(1) <= outputs_140108714735320(0);
        outputs_full_140108714735320(0) <= fifo_full_140108714735376(1);
        
        fifo_inputs_140108714735264(0) <= outputs_140108714735320(1);
        outputs_full_140108714735320(1) <= fifo_full_140108714735264(0);
        
        fifo_inputs_140108714735768(3) <= outputs_140108714735320(2);
        outputs_full_140108714735320(2) <= fifo_full_140108714735768(3);
        
        fifo_inputs_140108714734872(2) <= outputs_140108714735320(3);
        outputs_full_140108714735320(3) <= fifo_full_140108714734872(2);
        
        fifo_inputs_140108714735432(1) <= outputs_140108714735376(0);
        outputs_full_140108714735376(0) <= fifo_full_140108714735432(1);
        
        fifo_inputs_140108714735320(0) <= outputs_140108714735376(1);
        outputs_full_140108714735376(1) <= fifo_full_140108714735320(0);
        
        fifo_inputs_140108714735824(3) <= outputs_140108714735376(2);
        outputs_full_140108714735376(2) <= fifo_full_140108714735824(3);
        
        fifo_inputs_140108714734928(2) <= outputs_140108714735376(3);
        outputs_full_140108714735376(3) <= fifo_full_140108714734928(2);
        
        fifo_inputs_140108714735488(1) <= outputs_140108714735432(0);
        outputs_full_140108714735432(0) <= fifo_full_140108714735488(1);
        
        fifo_inputs_140108714735376(0) <= outputs_140108714735432(1);
        outputs_full_140108714735432(1) <= fifo_full_140108714735376(0);
        
        fifo_inputs_140108714735880(3) <= outputs_140108714735432(2);
        outputs_full_140108714735432(2) <= fifo_full_140108714735880(3);
        
        fifo_inputs_140108714734984(2) <= outputs_140108714735432(3);
        outputs_full_140108714735432(3) <= fifo_full_140108714734984(2);
        
        fifo_inputs_140108714735544(1) <= outputs_140108714735488(0);
        outputs_full_140108714735488(0) <= fifo_full_140108714735544(1);
        
        fifo_inputs_140108714735432(0) <= outputs_140108714735488(1);
        outputs_full_140108714735488(1) <= fifo_full_140108714735432(0);
        
        fifo_inputs_140108714735936(3) <= outputs_140108714735488(2);
        outputs_full_140108714735488(2) <= fifo_full_140108714735936(3);
        
        fifo_inputs_140108714735040(2) <= outputs_140108714735488(3);
        outputs_full_140108714735488(3) <= fifo_full_140108714735040(2);
        
        fifo_inputs_140108714735488(0) <= outputs_140108714735544(1);
        outputs_full_140108714735544(1) <= fifo_full_140108714735488(0);
        
        fifo_inputs_140108714735992(3) <= outputs_140108714735544(2);
        outputs_full_140108714735544(2) <= fifo_full_140108714735992(3);
        
        fifo_inputs_140108714735096(2) <= outputs_140108714735544(3);
        outputs_full_140108714735544(3) <= fifo_full_140108714735096(2);
        
        fifo_inputs_140108714735656(1) <= outputs_140108714735600(0);
        outputs_full_140108714735600(0) <= fifo_full_140108714735656(1);
        
        fifo_inputs_140108714736048(3) <= outputs_140108714735600(2);
        outputs_full_140108714735600(2) <= fifo_full_140108714736048(3);
        
        fifo_inputs_140108714735152(2) <= outputs_140108714735600(3);
        outputs_full_140108714735600(3) <= fifo_full_140108714735152(2);
        
        fifo_inputs_140108714735712(1) <= outputs_140108714735656(0);
        outputs_full_140108714735656(0) <= fifo_full_140108714735712(1);
        
        fifo_inputs_140108714735600(0) <= outputs_140108714735656(1);
        outputs_full_140108714735656(1) <= fifo_full_140108714735600(0);
        
        fifo_inputs_140108714736104(3) <= outputs_140108714735656(2);
        outputs_full_140108714735656(2) <= fifo_full_140108714736104(3);
        
        fifo_inputs_140108714735208(2) <= outputs_140108714735656(3);
        outputs_full_140108714735656(3) <= fifo_full_140108714735208(2);
        
        fifo_inputs_140108714735768(1) <= outputs_140108714735712(0);
        outputs_full_140108714735712(0) <= fifo_full_140108714735768(1);
        
        fifo_inputs_140108714735656(0) <= outputs_140108714735712(1);
        outputs_full_140108714735712(1) <= fifo_full_140108714735656(0);
        
        fifo_inputs_140108714736160(3) <= outputs_140108714735712(2);
        outputs_full_140108714735712(2) <= fifo_full_140108714736160(3);
        
        fifo_inputs_140108714735264(2) <= outputs_140108714735712(3);
        outputs_full_140108714735712(3) <= fifo_full_140108714735264(2);
        
        fifo_inputs_140108714735824(1) <= outputs_140108714735768(0);
        outputs_full_140108714735768(0) <= fifo_full_140108714735824(1);
        
        fifo_inputs_140108714735712(0) <= outputs_140108714735768(1);
        outputs_full_140108714735768(1) <= fifo_full_140108714735712(0);
        
        fifo_inputs_140108714736216(3) <= outputs_140108714735768(2);
        outputs_full_140108714735768(2) <= fifo_full_140108714736216(3);
        
        fifo_inputs_140108714735320(2) <= outputs_140108714735768(3);
        outputs_full_140108714735768(3) <= fifo_full_140108714735320(2);
        
        fifo_inputs_140108714735880(1) <= outputs_140108714735824(0);
        outputs_full_140108714735824(0) <= fifo_full_140108714735880(1);
        
        fifo_inputs_140108714735768(0) <= outputs_140108714735824(1);
        outputs_full_140108714735824(1) <= fifo_full_140108714735768(0);
        
        fifo_inputs_140108714736272(3) <= outputs_140108714735824(2);
        outputs_full_140108714735824(2) <= fifo_full_140108714736272(3);
        
        fifo_inputs_140108714735376(2) <= outputs_140108714735824(3);
        outputs_full_140108714735824(3) <= fifo_full_140108714735376(2);
        
        fifo_inputs_140108714735936(1) <= outputs_140108714735880(0);
        outputs_full_140108714735880(0) <= fifo_full_140108714735936(1);
        
        fifo_inputs_140108714735824(0) <= outputs_140108714735880(1);
        outputs_full_140108714735880(1) <= fifo_full_140108714735824(0);
        
        fifo_inputs_140108714736328(3) <= outputs_140108714735880(2);
        outputs_full_140108714735880(2) <= fifo_full_140108714736328(3);
        
        fifo_inputs_140108714735432(2) <= outputs_140108714735880(3);
        outputs_full_140108714735880(3) <= fifo_full_140108714735432(2);
        
        fifo_inputs_140108714735992(1) <= outputs_140108714735936(0);
        outputs_full_140108714735936(0) <= fifo_full_140108714735992(1);
        
        fifo_inputs_140108714735880(0) <= outputs_140108714735936(1);
        outputs_full_140108714735936(1) <= fifo_full_140108714735880(0);
        
        fifo_inputs_140108714736384(3) <= outputs_140108714735936(2);
        outputs_full_140108714735936(2) <= fifo_full_140108714736384(3);
        
        fifo_inputs_140108714735488(2) <= outputs_140108714735936(3);
        outputs_full_140108714735936(3) <= fifo_full_140108714735488(2);
        
        fifo_inputs_140108714735936(0) <= outputs_140108714735992(1);
        outputs_full_140108714735992(1) <= fifo_full_140108714735936(0);
        
        fifo_inputs_140108714736440(3) <= outputs_140108714735992(2);
        outputs_full_140108714735992(2) <= fifo_full_140108714736440(3);
        
        fifo_inputs_140108714735544(2) <= outputs_140108714735992(3);
        outputs_full_140108714735992(3) <= fifo_full_140108714735544(2);
        
        fifo_inputs_140108714736104(1) <= outputs_140108714736048(0);
        outputs_full_140108714736048(0) <= fifo_full_140108714736104(1);
        
        fifo_inputs_140108714735600(2) <= outputs_140108714736048(3);
        outputs_full_140108714736048(3) <= fifo_full_140108714735600(2);
        
        fifo_inputs_140108714736160(1) <= outputs_140108714736104(0);
        outputs_full_140108714736104(0) <= fifo_full_140108714736160(1);
        
        fifo_inputs_140108714736048(0) <= outputs_140108714736104(1);
        outputs_full_140108714736104(1) <= fifo_full_140108714736048(0);
        
        fifo_inputs_140108714735656(2) <= outputs_140108714736104(3);
        outputs_full_140108714736104(3) <= fifo_full_140108714735656(2);
        
        fifo_inputs_140108714736216(1) <= outputs_140108714736160(0);
        outputs_full_140108714736160(0) <= fifo_full_140108714736216(1);
        
        fifo_inputs_140108714736104(0) <= outputs_140108714736160(1);
        outputs_full_140108714736160(1) <= fifo_full_140108714736104(0);
        
        fifo_inputs_140108714735712(2) <= outputs_140108714736160(3);
        outputs_full_140108714736160(3) <= fifo_full_140108714735712(2);
        
        fifo_inputs_140108714736272(1) <= outputs_140108714736216(0);
        outputs_full_140108714736216(0) <= fifo_full_140108714736272(1);
        
        fifo_inputs_140108714736160(0) <= outputs_140108714736216(1);
        outputs_full_140108714736216(1) <= fifo_full_140108714736160(0);
        
        fifo_inputs_140108714735768(2) <= outputs_140108714736216(3);
        outputs_full_140108714736216(3) <= fifo_full_140108714735768(2);
        
        fifo_inputs_140108714736328(1) <= outputs_140108714736272(0);
        outputs_full_140108714736272(0) <= fifo_full_140108714736328(1);
        
        fifo_inputs_140108714736216(0) <= outputs_140108714736272(1);
        outputs_full_140108714736272(1) <= fifo_full_140108714736216(0);
        
        fifo_inputs_140108714735824(2) <= outputs_140108714736272(3);
        outputs_full_140108714736272(3) <= fifo_full_140108714735824(2);
        
        fifo_inputs_140108714736384(1) <= outputs_140108714736328(0);
        outputs_full_140108714736328(0) <= fifo_full_140108714736384(1);
        
        fifo_inputs_140108714736272(0) <= outputs_140108714736328(1);
        outputs_full_140108714736328(1) <= fifo_full_140108714736272(0);
        
        fifo_inputs_140108714735880(2) <= outputs_140108714736328(3);
        outputs_full_140108714736328(3) <= fifo_full_140108714735880(2);
        
        fifo_inputs_140108714736440(1) <= outputs_140108714736384(0);
        outputs_full_140108714736384(0) <= fifo_full_140108714736440(1);
        
        fifo_inputs_140108714736328(0) <= outputs_140108714736384(1);
        outputs_full_140108714736384(1) <= fifo_full_140108714736328(0);
        
        fifo_inputs_140108714735936(2) <= outputs_140108714736384(3);
        outputs_full_140108714736384(3) <= fifo_full_140108714735936(2);
        
        fifo_inputs_140108714736384(0) <= outputs_140108714736440(1);
        outputs_full_140108714736440(1) <= fifo_full_140108714736384(0);
        
        fifo_inputs_140108714735992(2) <= outputs_140108714736440(3);
        outputs_full_140108714736440(3) <= fifo_full_140108714735992(2);
        

    
        core_inst_140108714687736: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714687736,
            fifo_full => fifo_full_140108714687736,
            outputs => outputs_140108714687736,
            outputs_full => outputs_full_140108714687736
        );
        
        core_inst_140108714687960: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714687960,
            fifo_full => fifo_full_140108714687960,
            outputs => outputs_140108714687960,
            outputs_full => outputs_full_140108714687960
        );
        
        core_inst_140108714687904: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714687904,
            fifo_full => fifo_full_140108714687904,
            outputs => outputs_140108714687904,
            outputs_full => outputs_full_140108714687904
        );
        
        core_inst_140108714688016: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714688016,
            fifo_full => fifo_full_140108714688016,
            outputs => outputs_140108714688016,
            outputs_full => outputs_full_140108714688016
        );
        
        core_inst_140108714688072: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714688072,
            fifo_full => fifo_full_140108714688072,
            outputs => outputs_140108714688072,
            outputs_full => outputs_full_140108714688072
        );
        
        core_inst_140108714688128: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714688128,
            fifo_full => fifo_full_140108714688128,
            outputs => outputs_140108714688128,
            outputs_full => outputs_full_140108714688128
        );
        
        core_inst_140108714688184: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714688184,
            fifo_full => fifo_full_140108714688184,
            outputs => outputs_140108714688184,
            outputs_full => outputs_full_140108714688184
        );
        
        core_inst_140108714688240: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714688240,
            fifo_full => fifo_full_140108714688240,
            outputs => outputs_140108714688240,
            outputs_full => outputs_full_140108714688240
        );
        
        core_inst_140108714688296: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714688296,
            fifo_full => fifo_full_140108714688296,
            outputs => outputs_140108714688296,
            outputs_full => outputs_full_140108714688296
        );
        
        core_inst_140108714687848: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714687848,
            fifo_full => fifo_full_140108714687848,
            outputs => outputs_140108714687848,
            outputs_full => outputs_full_140108714687848
        );
        
        core_inst_140108714688352: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714688352,
            fifo_full => fifo_full_140108714688352,
            outputs => outputs_140108714688352,
            outputs_full => outputs_full_140108714688352
        );
        
        core_inst_140108714688408: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714688408,
            fifo_full => fifo_full_140108714688408,
            outputs => outputs_140108714688408,
            outputs_full => outputs_full_140108714688408
        );
        
        core_inst_140108714688464: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714688464,
            fifo_full => fifo_full_140108714688464,
            outputs => outputs_140108714688464,
            outputs_full => outputs_full_140108714688464
        );
        
        core_inst_140108714733640: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714733640,
            fifo_full => fifo_full_140108714733640,
            outputs => outputs_140108714733640,
            outputs_full => outputs_full_140108714733640
        );
        
        core_inst_140108714733696: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714733696,
            fifo_full => fifo_full_140108714733696,
            outputs => outputs_140108714733696,
            outputs_full => outputs_full_140108714733696
        );
        
        core_inst_140108714733752: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714733752,
            fifo_full => fifo_full_140108714733752,
            outputs => outputs_140108714733752,
            outputs_full => outputs_full_140108714733752
        );
        
        core_inst_140108714733808: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714733808,
            fifo_full => fifo_full_140108714733808,
            outputs => outputs_140108714733808,
            outputs_full => outputs_full_140108714733808
        );
        
        core_inst_140108714733864: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714733864,
            fifo_full => fifo_full_140108714733864,
            outputs => outputs_140108714733864,
            outputs_full => outputs_full_140108714733864
        );
        
        core_inst_140108714733920: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714733920,
            fifo_full => fifo_full_140108714733920,
            outputs => outputs_140108714733920,
            outputs_full => outputs_full_140108714733920
        );
        
        core_inst_140108714733976: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714733976,
            fifo_full => fifo_full_140108714733976,
            outputs => outputs_140108714733976,
            outputs_full => outputs_full_140108714733976
        );
        
        core_inst_140108714734032: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714734032,
            fifo_full => fifo_full_140108714734032,
            outputs => outputs_140108714734032,
            outputs_full => outputs_full_140108714734032
        );
        
        core_inst_140108714734088: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714734088,
            fifo_full => fifo_full_140108714734088,
            outputs => outputs_140108714734088,
            outputs_full => outputs_full_140108714734088
        );
        
        core_inst_140108714734144: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714734144,
            fifo_full => fifo_full_140108714734144,
            outputs => outputs_140108714734144,
            outputs_full => outputs_full_140108714734144
        );
        
        core_inst_140108714734200: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714734200,
            fifo_full => fifo_full_140108714734200,
            outputs => outputs_140108714734200,
            outputs_full => outputs_full_140108714734200
        );
        
        core_inst_140108714734256: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714734256,
            fifo_full => fifo_full_140108714734256,
            outputs => outputs_140108714734256,
            outputs_full => outputs_full_140108714734256
        );
        
        core_inst_140108714734312: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714734312,
            fifo_full => fifo_full_140108714734312,
            outputs => outputs_140108714734312,
            outputs_full => outputs_full_140108714734312
        );
        
        core_inst_140108714734368: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714734368,
            fifo_full => fifo_full_140108714734368,
            outputs => outputs_140108714734368,
            outputs_full => outputs_full_140108714734368
        );
        
        core_inst_140108714734424: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714734424,
            fifo_full => fifo_full_140108714734424,
            outputs => outputs_140108714734424,
            outputs_full => outputs_full_140108714734424
        );
        
        core_inst_140108714734480: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714734480,
            fifo_full => fifo_full_140108714734480,
            outputs => outputs_140108714734480,
            outputs_full => outputs_full_140108714734480
        );
        
        core_inst_140108714734536: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714734536,
            fifo_full => fifo_full_140108714734536,
            outputs => outputs_140108714734536,
            outputs_full => outputs_full_140108714734536
        );
        
        core_inst_140108714734592: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714734592,
            fifo_full => fifo_full_140108714734592,
            outputs => outputs_140108714734592,
            outputs_full => outputs_full_140108714734592
        );
        
        core_inst_140108714734648: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714734648,
            fifo_full => fifo_full_140108714734648,
            outputs => outputs_140108714734648,
            outputs_full => outputs_full_140108714734648
        );
        
        core_inst_140108714734704: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714734704,
            fifo_full => fifo_full_140108714734704,
            outputs => outputs_140108714734704,
            outputs_full => outputs_full_140108714734704
        );
        
        core_inst_140108714734760: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714734760,
            fifo_full => fifo_full_140108714734760,
            outputs => outputs_140108714734760,
            outputs_full => outputs_full_140108714734760
        );
        
        core_inst_140108714734816: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714734816,
            fifo_full => fifo_full_140108714734816,
            outputs => outputs_140108714734816,
            outputs_full => outputs_full_140108714734816
        );
        
        core_inst_140108714734872: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714734872,
            fifo_full => fifo_full_140108714734872,
            outputs => outputs_140108714734872,
            outputs_full => outputs_full_140108714734872
        );
        
        core_inst_140108714734928: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714734928,
            fifo_full => fifo_full_140108714734928,
            outputs => outputs_140108714734928,
            outputs_full => outputs_full_140108714734928
        );
        
        core_inst_140108714734984: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714734984,
            fifo_full => fifo_full_140108714734984,
            outputs => outputs_140108714734984,
            outputs_full => outputs_full_140108714734984
        );
        
        core_inst_140108714735040: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714735040,
            fifo_full => fifo_full_140108714735040,
            outputs => outputs_140108714735040,
            outputs_full => outputs_full_140108714735040
        );
        
        core_inst_140108714735096: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714735096,
            fifo_full => fifo_full_140108714735096,
            outputs => outputs_140108714735096,
            outputs_full => outputs_full_140108714735096
        );
        
        core_inst_140108714735152: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714735152,
            fifo_full => fifo_full_140108714735152,
            outputs => outputs_140108714735152,
            outputs_full => outputs_full_140108714735152
        );
        
        core_inst_140108714735208: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714735208,
            fifo_full => fifo_full_140108714735208,
            outputs => outputs_140108714735208,
            outputs_full => outputs_full_140108714735208
        );
        
        core_inst_140108714735264: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714735264,
            fifo_full => fifo_full_140108714735264,
            outputs => outputs_140108714735264,
            outputs_full => outputs_full_140108714735264
        );
        
        core_inst_140108714735320: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714735320,
            fifo_full => fifo_full_140108714735320,
            outputs => outputs_140108714735320,
            outputs_full => outputs_full_140108714735320
        );
        
        core_inst_140108714735376: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714735376,
            fifo_full => fifo_full_140108714735376,
            outputs => outputs_140108714735376,
            outputs_full => outputs_full_140108714735376
        );
        
        core_inst_140108714735432: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714735432,
            fifo_full => fifo_full_140108714735432,
            outputs => outputs_140108714735432,
            outputs_full => outputs_full_140108714735432
        );
        
        core_inst_140108714735488: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714735488,
            fifo_full => fifo_full_140108714735488,
            outputs => outputs_140108714735488,
            outputs_full => outputs_full_140108714735488
        );
        
        core_inst_140108714735544: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714735544,
            fifo_full => fifo_full_140108714735544,
            outputs => outputs_140108714735544,
            outputs_full => outputs_full_140108714735544
        );
        
        core_inst_140108714735600: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714735600,
            fifo_full => fifo_full_140108714735600,
            outputs => outputs_140108714735600,
            outputs_full => outputs_full_140108714735600
        );
        
        core_inst_140108714735656: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714735656,
            fifo_full => fifo_full_140108714735656,
            outputs => outputs_140108714735656,
            outputs_full => outputs_full_140108714735656
        );
        
        core_inst_140108714735712: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714735712,
            fifo_full => fifo_full_140108714735712,
            outputs => outputs_140108714735712,
            outputs_full => outputs_full_140108714735712
        );
        
        core_inst_140108714735768: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714735768,
            fifo_full => fifo_full_140108714735768,
            outputs => outputs_140108714735768,
            outputs_full => outputs_full_140108714735768
        );
        
        core_inst_140108714735824: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714735824,
            fifo_full => fifo_full_140108714735824,
            outputs => outputs_140108714735824,
            outputs_full => outputs_full_140108714735824
        );
        
        core_inst_140108714735880: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714735880,
            fifo_full => fifo_full_140108714735880,
            outputs => outputs_140108714735880,
            outputs_full => outputs_full_140108714735880
        );
        
        core_inst_140108714735936: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714735936,
            fifo_full => fifo_full_140108714735936,
            outputs => outputs_140108714735936,
            outputs_full => outputs_full_140108714735936
        );
        
        core_inst_140108714735992: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714735992,
            fifo_full => fifo_full_140108714735992,
            outputs => outputs_140108714735992,
            outputs_full => outputs_full_140108714735992
        );
        
        core_inst_140108714736048: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714736048,
            fifo_full => fifo_full_140108714736048,
            outputs => outputs_140108714736048,
            outputs_full => outputs_full_140108714736048
        );
        
        core_inst_140108714736104: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714736104,
            fifo_full => fifo_full_140108714736104,
            outputs => outputs_140108714736104,
            outputs_full => outputs_full_140108714736104
        );
        
        core_inst_140108714736160: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714736160,
            fifo_full => fifo_full_140108714736160,
            outputs => outputs_140108714736160,
            outputs_full => outputs_full_140108714736160
        );
        
        core_inst_140108714736216: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714736216,
            fifo_full => fifo_full_140108714736216,
            outputs => outputs_140108714736216,
            outputs_full => outputs_full_140108714736216
        );
        
        core_inst_140108714736272: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714736272,
            fifo_full => fifo_full_140108714736272,
            outputs => outputs_140108714736272,
            outputs_full => outputs_full_140108714736272
        );
        
        core_inst_140108714736328: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714736328,
            fifo_full => fifo_full_140108714736328,
            outputs => outputs_140108714736328,
            outputs_full => outputs_full_140108714736328
        );
        
        core_inst_140108714736384: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714736384,
            fifo_full => fifo_full_140108714736384,
            outputs => outputs_140108714736384,
            outputs_full => outputs_full_140108714736384
        );
        
        core_inst_140108714736440: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140108714736440,
            fifo_full => fifo_full_140108714736440,
            outputs => outputs_140108714736440,
            outputs_full => outputs_full_140108714736440
        );
        

end behav;

