
library ieee;
use ieee.std_logic_1164.all;
use work.core_config.all;
use work.all;

entity Bichain256 is
    port (
        clk: in std_logic;
        clk_en: in std_logic;
        reset: in std_logic;
        addr: in ram_addr;
        data: in word;
        we: in std_logic;
        fifo_inputs: in core_fifo_inputs_t;
        fifo_full: out std_logic_vector(0 to NUM_CORE_FIFOS-1);
        outputs: out core_fifo_inputs_t;
        outputs_full: in std_logic_vector(0 to NUM_CORE_FIFOS-1)
    );
end Bichain256;

architecture behav of Bichain256 is

    
        signal fifo_inputs_140423305571464: core_fifo_inputs_t;
        signal fifo_full_140423305571464: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305571464: core_fifo_inputs_t;
        signal outputs_full_140423305571464: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305571408: core_fifo_inputs_t;
        signal fifo_full_140423305571408: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305571408: core_fifo_inputs_t;
        signal outputs_full_140423305571408: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305571632: core_fifo_inputs_t;
        signal fifo_full_140423305571632: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305571632: core_fifo_inputs_t;
        signal outputs_full_140423305571632: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305571688: core_fifo_inputs_t;
        signal fifo_full_140423305571688: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305571688: core_fifo_inputs_t;
        signal outputs_full_140423305571688: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305571744: core_fifo_inputs_t;
        signal fifo_full_140423305571744: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305571744: core_fifo_inputs_t;
        signal outputs_full_140423305571744: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305571576: core_fifo_inputs_t;
        signal fifo_full_140423305571576: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305571576: core_fifo_inputs_t;
        signal outputs_full_140423305571576: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305571800: core_fifo_inputs_t;
        signal fifo_full_140423305571800: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305571800: core_fifo_inputs_t;
        signal outputs_full_140423305571800: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305571856: core_fifo_inputs_t;
        signal fifo_full_140423305571856: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305571856: core_fifo_inputs_t;
        signal outputs_full_140423305571856: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305571912: core_fifo_inputs_t;
        signal fifo_full_140423305571912: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305571912: core_fifo_inputs_t;
        signal outputs_full_140423305571912: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305571968: core_fifo_inputs_t;
        signal fifo_full_140423305571968: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305571968: core_fifo_inputs_t;
        signal outputs_full_140423305571968: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305571520: core_fifo_inputs_t;
        signal fifo_full_140423305571520: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305571520: core_fifo_inputs_t;
        signal outputs_full_140423305571520: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305572024: core_fifo_inputs_t;
        signal fifo_full_140423305572024: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305572024: core_fifo_inputs_t;
        signal outputs_full_140423305572024: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305572080: core_fifo_inputs_t;
        signal fifo_full_140423305572080: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305572080: core_fifo_inputs_t;
        signal outputs_full_140423305572080: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305572136: core_fifo_inputs_t;
        signal fifo_full_140423305572136: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305572136: core_fifo_inputs_t;
        signal outputs_full_140423305572136: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305572192: core_fifo_inputs_t;
        signal fifo_full_140423305572192: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305572192: core_fifo_inputs_t;
        signal outputs_full_140423305572192: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305572248: core_fifo_inputs_t;
        signal fifo_full_140423305572248: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305572248: core_fifo_inputs_t;
        signal outputs_full_140423305572248: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305572304: core_fifo_inputs_t;
        signal fifo_full_140423305572304: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305572304: core_fifo_inputs_t;
        signal outputs_full_140423305572304: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305621576: core_fifo_inputs_t;
        signal fifo_full_140423305621576: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305621576: core_fifo_inputs_t;
        signal outputs_full_140423305621576: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305621632: core_fifo_inputs_t;
        signal fifo_full_140423305621632: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305621632: core_fifo_inputs_t;
        signal outputs_full_140423305621632: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305621688: core_fifo_inputs_t;
        signal fifo_full_140423305621688: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305621688: core_fifo_inputs_t;
        signal outputs_full_140423305621688: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305621744: core_fifo_inputs_t;
        signal fifo_full_140423305621744: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305621744: core_fifo_inputs_t;
        signal outputs_full_140423305621744: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305621800: core_fifo_inputs_t;
        signal fifo_full_140423305621800: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305621800: core_fifo_inputs_t;
        signal outputs_full_140423305621800: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305621856: core_fifo_inputs_t;
        signal fifo_full_140423305621856: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305621856: core_fifo_inputs_t;
        signal outputs_full_140423305621856: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305621912: core_fifo_inputs_t;
        signal fifo_full_140423305621912: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305621912: core_fifo_inputs_t;
        signal outputs_full_140423305621912: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305621968: core_fifo_inputs_t;
        signal fifo_full_140423305621968: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305621968: core_fifo_inputs_t;
        signal outputs_full_140423305621968: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305622024: core_fifo_inputs_t;
        signal fifo_full_140423305622024: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305622024: core_fifo_inputs_t;
        signal outputs_full_140423305622024: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305622080: core_fifo_inputs_t;
        signal fifo_full_140423305622080: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305622080: core_fifo_inputs_t;
        signal outputs_full_140423305622080: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305622136: core_fifo_inputs_t;
        signal fifo_full_140423305622136: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305622136: core_fifo_inputs_t;
        signal outputs_full_140423305622136: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305622192: core_fifo_inputs_t;
        signal fifo_full_140423305622192: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305622192: core_fifo_inputs_t;
        signal outputs_full_140423305622192: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305622248: core_fifo_inputs_t;
        signal fifo_full_140423305622248: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305622248: core_fifo_inputs_t;
        signal outputs_full_140423305622248: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305622304: core_fifo_inputs_t;
        signal fifo_full_140423305622304: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305622304: core_fifo_inputs_t;
        signal outputs_full_140423305622304: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305622360: core_fifo_inputs_t;
        signal fifo_full_140423305622360: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305622360: core_fifo_inputs_t;
        signal outputs_full_140423305622360: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305622416: core_fifo_inputs_t;
        signal fifo_full_140423305622416: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305622416: core_fifo_inputs_t;
        signal outputs_full_140423305622416: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305622472: core_fifo_inputs_t;
        signal fifo_full_140423305622472: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305622472: core_fifo_inputs_t;
        signal outputs_full_140423305622472: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305622528: core_fifo_inputs_t;
        signal fifo_full_140423305622528: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305622528: core_fifo_inputs_t;
        signal outputs_full_140423305622528: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305622584: core_fifo_inputs_t;
        signal fifo_full_140423305622584: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305622584: core_fifo_inputs_t;
        signal outputs_full_140423305622584: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305622640: core_fifo_inputs_t;
        signal fifo_full_140423305622640: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305622640: core_fifo_inputs_t;
        signal outputs_full_140423305622640: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305622696: core_fifo_inputs_t;
        signal fifo_full_140423305622696: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305622696: core_fifo_inputs_t;
        signal outputs_full_140423305622696: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305622752: core_fifo_inputs_t;
        signal fifo_full_140423305622752: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305622752: core_fifo_inputs_t;
        signal outputs_full_140423305622752: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305622808: core_fifo_inputs_t;
        signal fifo_full_140423305622808: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305622808: core_fifo_inputs_t;
        signal outputs_full_140423305622808: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305622864: core_fifo_inputs_t;
        signal fifo_full_140423305622864: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305622864: core_fifo_inputs_t;
        signal outputs_full_140423305622864: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305622920: core_fifo_inputs_t;
        signal fifo_full_140423305622920: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305622920: core_fifo_inputs_t;
        signal outputs_full_140423305622920: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305622976: core_fifo_inputs_t;
        signal fifo_full_140423305622976: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305622976: core_fifo_inputs_t;
        signal outputs_full_140423305622976: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305623032: core_fifo_inputs_t;
        signal fifo_full_140423305623032: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305623032: core_fifo_inputs_t;
        signal outputs_full_140423305623032: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305623088: core_fifo_inputs_t;
        signal fifo_full_140423305623088: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305623088: core_fifo_inputs_t;
        signal outputs_full_140423305623088: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305623144: core_fifo_inputs_t;
        signal fifo_full_140423305623144: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305623144: core_fifo_inputs_t;
        signal outputs_full_140423305623144: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305623200: core_fifo_inputs_t;
        signal fifo_full_140423305623200: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305623200: core_fifo_inputs_t;
        signal outputs_full_140423305623200: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305623256: core_fifo_inputs_t;
        signal fifo_full_140423305623256: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305623256: core_fifo_inputs_t;
        signal outputs_full_140423305623256: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305623312: core_fifo_inputs_t;
        signal fifo_full_140423305623312: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305623312: core_fifo_inputs_t;
        signal outputs_full_140423305623312: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305623368: core_fifo_inputs_t;
        signal fifo_full_140423305623368: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305623368: core_fifo_inputs_t;
        signal outputs_full_140423305623368: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305623424: core_fifo_inputs_t;
        signal fifo_full_140423305623424: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305623424: core_fifo_inputs_t;
        signal outputs_full_140423305623424: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305623480: core_fifo_inputs_t;
        signal fifo_full_140423305623480: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305623480: core_fifo_inputs_t;
        signal outputs_full_140423305623480: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305623536: core_fifo_inputs_t;
        signal fifo_full_140423305623536: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305623536: core_fifo_inputs_t;
        signal outputs_full_140423305623536: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305623592: core_fifo_inputs_t;
        signal fifo_full_140423305623592: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305623592: core_fifo_inputs_t;
        signal outputs_full_140423305623592: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305623648: core_fifo_inputs_t;
        signal fifo_full_140423305623648: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305623648: core_fifo_inputs_t;
        signal outputs_full_140423305623648: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305623704: core_fifo_inputs_t;
        signal fifo_full_140423305623704: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305623704: core_fifo_inputs_t;
        signal outputs_full_140423305623704: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305623760: core_fifo_inputs_t;
        signal fifo_full_140423305623760: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305623760: core_fifo_inputs_t;
        signal outputs_full_140423305623760: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305623816: core_fifo_inputs_t;
        signal fifo_full_140423305623816: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305623816: core_fifo_inputs_t;
        signal outputs_full_140423305623816: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305623872: core_fifo_inputs_t;
        signal fifo_full_140423305623872: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305623872: core_fifo_inputs_t;
        signal outputs_full_140423305623872: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305623928: core_fifo_inputs_t;
        signal fifo_full_140423305623928: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305623928: core_fifo_inputs_t;
        signal outputs_full_140423305623928: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305623984: core_fifo_inputs_t;
        signal fifo_full_140423305623984: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305623984: core_fifo_inputs_t;
        signal outputs_full_140423305623984: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305624040: core_fifo_inputs_t;
        signal fifo_full_140423305624040: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305624040: core_fifo_inputs_t;
        signal outputs_full_140423305624040: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305624096: core_fifo_inputs_t;
        signal fifo_full_140423305624096: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305624096: core_fifo_inputs_t;
        signal outputs_full_140423305624096: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305624152: core_fifo_inputs_t;
        signal fifo_full_140423305624152: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305624152: core_fifo_inputs_t;
        signal outputs_full_140423305624152: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305624208: core_fifo_inputs_t;
        signal fifo_full_140423305624208: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305624208: core_fifo_inputs_t;
        signal outputs_full_140423305624208: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305624264: core_fifo_inputs_t;
        signal fifo_full_140423305624264: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305624264: core_fifo_inputs_t;
        signal outputs_full_140423305624264: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305624320: core_fifo_inputs_t;
        signal fifo_full_140423305624320: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305624320: core_fifo_inputs_t;
        signal outputs_full_140423305624320: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305624376: core_fifo_inputs_t;
        signal fifo_full_140423305624376: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305624376: core_fifo_inputs_t;
        signal outputs_full_140423305624376: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305624432: core_fifo_inputs_t;
        signal fifo_full_140423305624432: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305624432: core_fifo_inputs_t;
        signal outputs_full_140423305624432: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305624488: core_fifo_inputs_t;
        signal fifo_full_140423305624488: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305624488: core_fifo_inputs_t;
        signal outputs_full_140423305624488: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305624544: core_fifo_inputs_t;
        signal fifo_full_140423305624544: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305624544: core_fifo_inputs_t;
        signal outputs_full_140423305624544: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305624600: core_fifo_inputs_t;
        signal fifo_full_140423305624600: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305624600: core_fifo_inputs_t;
        signal outputs_full_140423305624600: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305624656: core_fifo_inputs_t;
        signal fifo_full_140423305624656: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305624656: core_fifo_inputs_t;
        signal outputs_full_140423305624656: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305624712: core_fifo_inputs_t;
        signal fifo_full_140423305624712: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305624712: core_fifo_inputs_t;
        signal outputs_full_140423305624712: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305624768: core_fifo_inputs_t;
        signal fifo_full_140423305624768: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305624768: core_fifo_inputs_t;
        signal outputs_full_140423305624768: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305624824: core_fifo_inputs_t;
        signal fifo_full_140423305624824: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305624824: core_fifo_inputs_t;
        signal outputs_full_140423305624824: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305624880: core_fifo_inputs_t;
        signal fifo_full_140423305624880: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305624880: core_fifo_inputs_t;
        signal outputs_full_140423305624880: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305624936: core_fifo_inputs_t;
        signal fifo_full_140423305624936: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305624936: core_fifo_inputs_t;
        signal outputs_full_140423305624936: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305624992: core_fifo_inputs_t;
        signal fifo_full_140423305624992: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305624992: core_fifo_inputs_t;
        signal outputs_full_140423305624992: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305625048: core_fifo_inputs_t;
        signal fifo_full_140423305625048: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305625048: core_fifo_inputs_t;
        signal outputs_full_140423305625048: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305625104: core_fifo_inputs_t;
        signal fifo_full_140423305625104: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305625104: core_fifo_inputs_t;
        signal outputs_full_140423305625104: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305625160: core_fifo_inputs_t;
        signal fifo_full_140423305625160: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305625160: core_fifo_inputs_t;
        signal outputs_full_140423305625160: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305625216: core_fifo_inputs_t;
        signal fifo_full_140423305625216: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305625216: core_fifo_inputs_t;
        signal outputs_full_140423305625216: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305625272: core_fifo_inputs_t;
        signal fifo_full_140423305625272: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305625272: core_fifo_inputs_t;
        signal outputs_full_140423305625272: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305625328: core_fifo_inputs_t;
        signal fifo_full_140423305625328: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305625328: core_fifo_inputs_t;
        signal outputs_full_140423305625328: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305625384: core_fifo_inputs_t;
        signal fifo_full_140423305625384: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305625384: core_fifo_inputs_t;
        signal outputs_full_140423305625384: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305625440: core_fifo_inputs_t;
        signal fifo_full_140423305625440: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305625440: core_fifo_inputs_t;
        signal outputs_full_140423305625440: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305625496: core_fifo_inputs_t;
        signal fifo_full_140423305625496: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305625496: core_fifo_inputs_t;
        signal outputs_full_140423305625496: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305625552: core_fifo_inputs_t;
        signal fifo_full_140423305625552: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305625552: core_fifo_inputs_t;
        signal outputs_full_140423305625552: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305642056: core_fifo_inputs_t;
        signal fifo_full_140423305642056: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305642056: core_fifo_inputs_t;
        signal outputs_full_140423305642056: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305642112: core_fifo_inputs_t;
        signal fifo_full_140423305642112: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305642112: core_fifo_inputs_t;
        signal outputs_full_140423305642112: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305642168: core_fifo_inputs_t;
        signal fifo_full_140423305642168: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305642168: core_fifo_inputs_t;
        signal outputs_full_140423305642168: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305642224: core_fifo_inputs_t;
        signal fifo_full_140423305642224: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305642224: core_fifo_inputs_t;
        signal outputs_full_140423305642224: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305642280: core_fifo_inputs_t;
        signal fifo_full_140423305642280: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305642280: core_fifo_inputs_t;
        signal outputs_full_140423305642280: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305642336: core_fifo_inputs_t;
        signal fifo_full_140423305642336: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305642336: core_fifo_inputs_t;
        signal outputs_full_140423305642336: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305642392: core_fifo_inputs_t;
        signal fifo_full_140423305642392: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305642392: core_fifo_inputs_t;
        signal outputs_full_140423305642392: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305642448: core_fifo_inputs_t;
        signal fifo_full_140423305642448: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305642448: core_fifo_inputs_t;
        signal outputs_full_140423305642448: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305642504: core_fifo_inputs_t;
        signal fifo_full_140423305642504: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305642504: core_fifo_inputs_t;
        signal outputs_full_140423305642504: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305642560: core_fifo_inputs_t;
        signal fifo_full_140423305642560: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305642560: core_fifo_inputs_t;
        signal outputs_full_140423305642560: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305642616: core_fifo_inputs_t;
        signal fifo_full_140423305642616: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305642616: core_fifo_inputs_t;
        signal outputs_full_140423305642616: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305642672: core_fifo_inputs_t;
        signal fifo_full_140423305642672: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305642672: core_fifo_inputs_t;
        signal outputs_full_140423305642672: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305642728: core_fifo_inputs_t;
        signal fifo_full_140423305642728: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305642728: core_fifo_inputs_t;
        signal outputs_full_140423305642728: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305642784: core_fifo_inputs_t;
        signal fifo_full_140423305642784: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305642784: core_fifo_inputs_t;
        signal outputs_full_140423305642784: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305642840: core_fifo_inputs_t;
        signal fifo_full_140423305642840: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305642840: core_fifo_inputs_t;
        signal outputs_full_140423305642840: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305642896: core_fifo_inputs_t;
        signal fifo_full_140423305642896: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305642896: core_fifo_inputs_t;
        signal outputs_full_140423305642896: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305642952: core_fifo_inputs_t;
        signal fifo_full_140423305642952: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305642952: core_fifo_inputs_t;
        signal outputs_full_140423305642952: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305643008: core_fifo_inputs_t;
        signal fifo_full_140423305643008: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305643008: core_fifo_inputs_t;
        signal outputs_full_140423305643008: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305643064: core_fifo_inputs_t;
        signal fifo_full_140423305643064: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305643064: core_fifo_inputs_t;
        signal outputs_full_140423305643064: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305643120: core_fifo_inputs_t;
        signal fifo_full_140423305643120: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305643120: core_fifo_inputs_t;
        signal outputs_full_140423305643120: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305643176: core_fifo_inputs_t;
        signal fifo_full_140423305643176: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305643176: core_fifo_inputs_t;
        signal outputs_full_140423305643176: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305643232: core_fifo_inputs_t;
        signal fifo_full_140423305643232: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305643232: core_fifo_inputs_t;
        signal outputs_full_140423305643232: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305643288: core_fifo_inputs_t;
        signal fifo_full_140423305643288: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305643288: core_fifo_inputs_t;
        signal outputs_full_140423305643288: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305643344: core_fifo_inputs_t;
        signal fifo_full_140423305643344: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305643344: core_fifo_inputs_t;
        signal outputs_full_140423305643344: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305643400: core_fifo_inputs_t;
        signal fifo_full_140423305643400: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305643400: core_fifo_inputs_t;
        signal outputs_full_140423305643400: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305643456: core_fifo_inputs_t;
        signal fifo_full_140423305643456: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305643456: core_fifo_inputs_t;
        signal outputs_full_140423305643456: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305643512: core_fifo_inputs_t;
        signal fifo_full_140423305643512: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305643512: core_fifo_inputs_t;
        signal outputs_full_140423305643512: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305643568: core_fifo_inputs_t;
        signal fifo_full_140423305643568: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305643568: core_fifo_inputs_t;
        signal outputs_full_140423305643568: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305643624: core_fifo_inputs_t;
        signal fifo_full_140423305643624: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305643624: core_fifo_inputs_t;
        signal outputs_full_140423305643624: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305643680: core_fifo_inputs_t;
        signal fifo_full_140423305643680: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305643680: core_fifo_inputs_t;
        signal outputs_full_140423305643680: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305643736: core_fifo_inputs_t;
        signal fifo_full_140423305643736: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305643736: core_fifo_inputs_t;
        signal outputs_full_140423305643736: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305643792: core_fifo_inputs_t;
        signal fifo_full_140423305643792: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305643792: core_fifo_inputs_t;
        signal outputs_full_140423305643792: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305643848: core_fifo_inputs_t;
        signal fifo_full_140423305643848: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305643848: core_fifo_inputs_t;
        signal outputs_full_140423305643848: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305643904: core_fifo_inputs_t;
        signal fifo_full_140423305643904: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305643904: core_fifo_inputs_t;
        signal outputs_full_140423305643904: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305643960: core_fifo_inputs_t;
        signal fifo_full_140423305643960: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305643960: core_fifo_inputs_t;
        signal outputs_full_140423305643960: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305644016: core_fifo_inputs_t;
        signal fifo_full_140423305644016: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305644016: core_fifo_inputs_t;
        signal outputs_full_140423305644016: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305644072: core_fifo_inputs_t;
        signal fifo_full_140423305644072: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305644072: core_fifo_inputs_t;
        signal outputs_full_140423305644072: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305644128: core_fifo_inputs_t;
        signal fifo_full_140423305644128: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305644128: core_fifo_inputs_t;
        signal outputs_full_140423305644128: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305644184: core_fifo_inputs_t;
        signal fifo_full_140423305644184: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305644184: core_fifo_inputs_t;
        signal outputs_full_140423305644184: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305644240: core_fifo_inputs_t;
        signal fifo_full_140423305644240: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305644240: core_fifo_inputs_t;
        signal outputs_full_140423305644240: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305644296: core_fifo_inputs_t;
        signal fifo_full_140423305644296: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305644296: core_fifo_inputs_t;
        signal outputs_full_140423305644296: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305644352: core_fifo_inputs_t;
        signal fifo_full_140423305644352: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305644352: core_fifo_inputs_t;
        signal outputs_full_140423305644352: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305644408: core_fifo_inputs_t;
        signal fifo_full_140423305644408: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305644408: core_fifo_inputs_t;
        signal outputs_full_140423305644408: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305644464: core_fifo_inputs_t;
        signal fifo_full_140423305644464: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305644464: core_fifo_inputs_t;
        signal outputs_full_140423305644464: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305644520: core_fifo_inputs_t;
        signal fifo_full_140423305644520: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305644520: core_fifo_inputs_t;
        signal outputs_full_140423305644520: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305644576: core_fifo_inputs_t;
        signal fifo_full_140423305644576: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305644576: core_fifo_inputs_t;
        signal outputs_full_140423305644576: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305644632: core_fifo_inputs_t;
        signal fifo_full_140423305644632: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305644632: core_fifo_inputs_t;
        signal outputs_full_140423305644632: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305644688: core_fifo_inputs_t;
        signal fifo_full_140423305644688: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305644688: core_fifo_inputs_t;
        signal outputs_full_140423305644688: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305644744: core_fifo_inputs_t;
        signal fifo_full_140423305644744: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305644744: core_fifo_inputs_t;
        signal outputs_full_140423305644744: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305644800: core_fifo_inputs_t;
        signal fifo_full_140423305644800: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305644800: core_fifo_inputs_t;
        signal outputs_full_140423305644800: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305644856: core_fifo_inputs_t;
        signal fifo_full_140423305644856: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305644856: core_fifo_inputs_t;
        signal outputs_full_140423305644856: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305644912: core_fifo_inputs_t;
        signal fifo_full_140423305644912: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305644912: core_fifo_inputs_t;
        signal outputs_full_140423305644912: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305644968: core_fifo_inputs_t;
        signal fifo_full_140423305644968: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305644968: core_fifo_inputs_t;
        signal outputs_full_140423305644968: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305645024: core_fifo_inputs_t;
        signal fifo_full_140423305645024: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305645024: core_fifo_inputs_t;
        signal outputs_full_140423305645024: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305645080: core_fifo_inputs_t;
        signal fifo_full_140423305645080: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305645080: core_fifo_inputs_t;
        signal outputs_full_140423305645080: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305645136: core_fifo_inputs_t;
        signal fifo_full_140423305645136: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305645136: core_fifo_inputs_t;
        signal outputs_full_140423305645136: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305645192: core_fifo_inputs_t;
        signal fifo_full_140423305645192: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305645192: core_fifo_inputs_t;
        signal outputs_full_140423305645192: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305645248: core_fifo_inputs_t;
        signal fifo_full_140423305645248: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305645248: core_fifo_inputs_t;
        signal outputs_full_140423305645248: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305645304: core_fifo_inputs_t;
        signal fifo_full_140423305645304: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305645304: core_fifo_inputs_t;
        signal outputs_full_140423305645304: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305645360: core_fifo_inputs_t;
        signal fifo_full_140423305645360: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305645360: core_fifo_inputs_t;
        signal outputs_full_140423305645360: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305645416: core_fifo_inputs_t;
        signal fifo_full_140423305645416: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305645416: core_fifo_inputs_t;
        signal outputs_full_140423305645416: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305645472: core_fifo_inputs_t;
        signal fifo_full_140423305645472: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305645472: core_fifo_inputs_t;
        signal outputs_full_140423305645472: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305645528: core_fifo_inputs_t;
        signal fifo_full_140423305645528: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305645528: core_fifo_inputs_t;
        signal outputs_full_140423305645528: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305645584: core_fifo_inputs_t;
        signal fifo_full_140423305645584: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305645584: core_fifo_inputs_t;
        signal outputs_full_140423305645584: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305645640: core_fifo_inputs_t;
        signal fifo_full_140423305645640: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305645640: core_fifo_inputs_t;
        signal outputs_full_140423305645640: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423329706112: core_fifo_inputs_t;
        signal fifo_full_140423329706112: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423329706112: core_fifo_inputs_t;
        signal outputs_full_140423329706112: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305571240: core_fifo_inputs_t;
        signal fifo_full_140423305571240: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305571240: core_fifo_inputs_t;
        signal outputs_full_140423305571240: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305571016: core_fifo_inputs_t;
        signal fifo_full_140423305571016: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305571016: core_fifo_inputs_t;
        signal outputs_full_140423305571016: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305571296: core_fifo_inputs_t;
        signal fifo_full_140423305571296: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305571296: core_fifo_inputs_t;
        signal outputs_full_140423305571296: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305571072: core_fifo_inputs_t;
        signal fifo_full_140423305571072: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305571072: core_fifo_inputs_t;
        signal outputs_full_140423305571072: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305571128: core_fifo_inputs_t;
        signal fifo_full_140423305571128: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305571128: core_fifo_inputs_t;
        signal outputs_full_140423305571128: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305645696: core_fifo_inputs_t;
        signal fifo_full_140423305645696: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305645696: core_fifo_inputs_t;
        signal outputs_full_140423305645696: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305645752: core_fifo_inputs_t;
        signal fifo_full_140423305645752: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305645752: core_fifo_inputs_t;
        signal outputs_full_140423305645752: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305645808: core_fifo_inputs_t;
        signal fifo_full_140423305645808: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305645808: core_fifo_inputs_t;
        signal outputs_full_140423305645808: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305645864: core_fifo_inputs_t;
        signal fifo_full_140423305645864: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305645864: core_fifo_inputs_t;
        signal outputs_full_140423305645864: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305645920: core_fifo_inputs_t;
        signal fifo_full_140423305645920: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305645920: core_fifo_inputs_t;
        signal outputs_full_140423305645920: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305645976: core_fifo_inputs_t;
        signal fifo_full_140423305645976: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305645976: core_fifo_inputs_t;
        signal outputs_full_140423305645976: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305646032: core_fifo_inputs_t;
        signal fifo_full_140423305646032: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305646032: core_fifo_inputs_t;
        signal outputs_full_140423305646032: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305662536: core_fifo_inputs_t;
        signal fifo_full_140423305662536: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305662536: core_fifo_inputs_t;
        signal outputs_full_140423305662536: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305662592: core_fifo_inputs_t;
        signal fifo_full_140423305662592: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305662592: core_fifo_inputs_t;
        signal outputs_full_140423305662592: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305662648: core_fifo_inputs_t;
        signal fifo_full_140423305662648: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305662648: core_fifo_inputs_t;
        signal outputs_full_140423305662648: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305662704: core_fifo_inputs_t;
        signal fifo_full_140423305662704: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305662704: core_fifo_inputs_t;
        signal outputs_full_140423305662704: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305662760: core_fifo_inputs_t;
        signal fifo_full_140423305662760: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305662760: core_fifo_inputs_t;
        signal outputs_full_140423305662760: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305662816: core_fifo_inputs_t;
        signal fifo_full_140423305662816: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305662816: core_fifo_inputs_t;
        signal outputs_full_140423305662816: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305662872: core_fifo_inputs_t;
        signal fifo_full_140423305662872: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305662872: core_fifo_inputs_t;
        signal outputs_full_140423305662872: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305662928: core_fifo_inputs_t;
        signal fifo_full_140423305662928: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305662928: core_fifo_inputs_t;
        signal outputs_full_140423305662928: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305662984: core_fifo_inputs_t;
        signal fifo_full_140423305662984: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305662984: core_fifo_inputs_t;
        signal outputs_full_140423305662984: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305663040: core_fifo_inputs_t;
        signal fifo_full_140423305663040: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305663040: core_fifo_inputs_t;
        signal outputs_full_140423305663040: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305663096: core_fifo_inputs_t;
        signal fifo_full_140423305663096: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305663096: core_fifo_inputs_t;
        signal outputs_full_140423305663096: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305663152: core_fifo_inputs_t;
        signal fifo_full_140423305663152: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305663152: core_fifo_inputs_t;
        signal outputs_full_140423305663152: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305663208: core_fifo_inputs_t;
        signal fifo_full_140423305663208: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305663208: core_fifo_inputs_t;
        signal outputs_full_140423305663208: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305663264: core_fifo_inputs_t;
        signal fifo_full_140423305663264: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305663264: core_fifo_inputs_t;
        signal outputs_full_140423305663264: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305663320: core_fifo_inputs_t;
        signal fifo_full_140423305663320: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305663320: core_fifo_inputs_t;
        signal outputs_full_140423305663320: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305663376: core_fifo_inputs_t;
        signal fifo_full_140423305663376: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305663376: core_fifo_inputs_t;
        signal outputs_full_140423305663376: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305663432: core_fifo_inputs_t;
        signal fifo_full_140423305663432: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305663432: core_fifo_inputs_t;
        signal outputs_full_140423305663432: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305663488: core_fifo_inputs_t;
        signal fifo_full_140423305663488: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305663488: core_fifo_inputs_t;
        signal outputs_full_140423305663488: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305663544: core_fifo_inputs_t;
        signal fifo_full_140423305663544: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305663544: core_fifo_inputs_t;
        signal outputs_full_140423305663544: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305663600: core_fifo_inputs_t;
        signal fifo_full_140423305663600: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305663600: core_fifo_inputs_t;
        signal outputs_full_140423305663600: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305663656: core_fifo_inputs_t;
        signal fifo_full_140423305663656: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305663656: core_fifo_inputs_t;
        signal outputs_full_140423305663656: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305663712: core_fifo_inputs_t;
        signal fifo_full_140423305663712: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305663712: core_fifo_inputs_t;
        signal outputs_full_140423305663712: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305663768: core_fifo_inputs_t;
        signal fifo_full_140423305663768: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305663768: core_fifo_inputs_t;
        signal outputs_full_140423305663768: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305663824: core_fifo_inputs_t;
        signal fifo_full_140423305663824: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305663824: core_fifo_inputs_t;
        signal outputs_full_140423305663824: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305663880: core_fifo_inputs_t;
        signal fifo_full_140423305663880: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305663880: core_fifo_inputs_t;
        signal outputs_full_140423305663880: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305663936: core_fifo_inputs_t;
        signal fifo_full_140423305663936: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305663936: core_fifo_inputs_t;
        signal outputs_full_140423305663936: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305663992: core_fifo_inputs_t;
        signal fifo_full_140423305663992: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305663992: core_fifo_inputs_t;
        signal outputs_full_140423305663992: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305664048: core_fifo_inputs_t;
        signal fifo_full_140423305664048: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305664048: core_fifo_inputs_t;
        signal outputs_full_140423305664048: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305664104: core_fifo_inputs_t;
        signal fifo_full_140423305664104: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305664104: core_fifo_inputs_t;
        signal outputs_full_140423305664104: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305664160: core_fifo_inputs_t;
        signal fifo_full_140423305664160: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305664160: core_fifo_inputs_t;
        signal outputs_full_140423305664160: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305664216: core_fifo_inputs_t;
        signal fifo_full_140423305664216: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305664216: core_fifo_inputs_t;
        signal outputs_full_140423305664216: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305664272: core_fifo_inputs_t;
        signal fifo_full_140423305664272: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305664272: core_fifo_inputs_t;
        signal outputs_full_140423305664272: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305664328: core_fifo_inputs_t;
        signal fifo_full_140423305664328: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305664328: core_fifo_inputs_t;
        signal outputs_full_140423305664328: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305664384: core_fifo_inputs_t;
        signal fifo_full_140423305664384: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305664384: core_fifo_inputs_t;
        signal outputs_full_140423305664384: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305664440: core_fifo_inputs_t;
        signal fifo_full_140423305664440: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305664440: core_fifo_inputs_t;
        signal outputs_full_140423305664440: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305664496: core_fifo_inputs_t;
        signal fifo_full_140423305664496: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305664496: core_fifo_inputs_t;
        signal outputs_full_140423305664496: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305664552: core_fifo_inputs_t;
        signal fifo_full_140423305664552: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305664552: core_fifo_inputs_t;
        signal outputs_full_140423305664552: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305664608: core_fifo_inputs_t;
        signal fifo_full_140423305664608: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305664608: core_fifo_inputs_t;
        signal outputs_full_140423305664608: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305664664: core_fifo_inputs_t;
        signal fifo_full_140423305664664: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305664664: core_fifo_inputs_t;
        signal outputs_full_140423305664664: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305664720: core_fifo_inputs_t;
        signal fifo_full_140423305664720: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305664720: core_fifo_inputs_t;
        signal outputs_full_140423305664720: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305664776: core_fifo_inputs_t;
        signal fifo_full_140423305664776: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305664776: core_fifo_inputs_t;
        signal outputs_full_140423305664776: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305664832: core_fifo_inputs_t;
        signal fifo_full_140423305664832: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305664832: core_fifo_inputs_t;
        signal outputs_full_140423305664832: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305664888: core_fifo_inputs_t;
        signal fifo_full_140423305664888: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305664888: core_fifo_inputs_t;
        signal outputs_full_140423305664888: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305664944: core_fifo_inputs_t;
        signal fifo_full_140423305664944: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305664944: core_fifo_inputs_t;
        signal outputs_full_140423305664944: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305665000: core_fifo_inputs_t;
        signal fifo_full_140423305665000: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305665000: core_fifo_inputs_t;
        signal outputs_full_140423305665000: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305665056: core_fifo_inputs_t;
        signal fifo_full_140423305665056: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305665056: core_fifo_inputs_t;
        signal outputs_full_140423305665056: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305665112: core_fifo_inputs_t;
        signal fifo_full_140423305665112: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305665112: core_fifo_inputs_t;
        signal outputs_full_140423305665112: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305665168: core_fifo_inputs_t;
        signal fifo_full_140423305665168: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305665168: core_fifo_inputs_t;
        signal outputs_full_140423305665168: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305665224: core_fifo_inputs_t;
        signal fifo_full_140423305665224: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305665224: core_fifo_inputs_t;
        signal outputs_full_140423305665224: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305665280: core_fifo_inputs_t;
        signal fifo_full_140423305665280: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305665280: core_fifo_inputs_t;
        signal outputs_full_140423305665280: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305665336: core_fifo_inputs_t;
        signal fifo_full_140423305665336: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305665336: core_fifo_inputs_t;
        signal outputs_full_140423305665336: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305665392: core_fifo_inputs_t;
        signal fifo_full_140423305665392: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305665392: core_fifo_inputs_t;
        signal outputs_full_140423305665392: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305665448: core_fifo_inputs_t;
        signal fifo_full_140423305665448: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305665448: core_fifo_inputs_t;
        signal outputs_full_140423305665448: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305665504: core_fifo_inputs_t;
        signal fifo_full_140423305665504: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305665504: core_fifo_inputs_t;
        signal outputs_full_140423305665504: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305665560: core_fifo_inputs_t;
        signal fifo_full_140423305665560: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305665560: core_fifo_inputs_t;
        signal outputs_full_140423305665560: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305665616: core_fifo_inputs_t;
        signal fifo_full_140423305665616: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305665616: core_fifo_inputs_t;
        signal outputs_full_140423305665616: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305665672: core_fifo_inputs_t;
        signal fifo_full_140423305665672: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305665672: core_fifo_inputs_t;
        signal outputs_full_140423305665672: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305665728: core_fifo_inputs_t;
        signal fifo_full_140423305665728: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305665728: core_fifo_inputs_t;
        signal outputs_full_140423305665728: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305665784: core_fifo_inputs_t;
        signal fifo_full_140423305665784: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305665784: core_fifo_inputs_t;
        signal outputs_full_140423305665784: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305665840: core_fifo_inputs_t;
        signal fifo_full_140423305665840: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305665840: core_fifo_inputs_t;
        signal outputs_full_140423305665840: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305665896: core_fifo_inputs_t;
        signal fifo_full_140423305665896: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305665896: core_fifo_inputs_t;
        signal outputs_full_140423305665896: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305665952: core_fifo_inputs_t;
        signal fifo_full_140423305665952: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305665952: core_fifo_inputs_t;
        signal outputs_full_140423305665952: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305666008: core_fifo_inputs_t;
        signal fifo_full_140423305666008: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305666008: core_fifo_inputs_t;
        signal outputs_full_140423305666008: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305666064: core_fifo_inputs_t;
        signal fifo_full_140423305666064: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305666064: core_fifo_inputs_t;
        signal outputs_full_140423305666064: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305666120: core_fifo_inputs_t;
        signal fifo_full_140423305666120: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305666120: core_fifo_inputs_t;
        signal outputs_full_140423305666120: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305666176: core_fifo_inputs_t;
        signal fifo_full_140423305666176: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305666176: core_fifo_inputs_t;
        signal outputs_full_140423305666176: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305666232: core_fifo_inputs_t;
        signal fifo_full_140423305666232: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305666232: core_fifo_inputs_t;
        signal outputs_full_140423305666232: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305666288: core_fifo_inputs_t;
        signal fifo_full_140423305666288: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305666288: core_fifo_inputs_t;
        signal outputs_full_140423305666288: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305666344: core_fifo_inputs_t;
        signal fifo_full_140423305666344: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305666344: core_fifo_inputs_t;
        signal outputs_full_140423305666344: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305666400: core_fifo_inputs_t;
        signal fifo_full_140423305666400: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305666400: core_fifo_inputs_t;
        signal outputs_full_140423305666400: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305666456: core_fifo_inputs_t;
        signal fifo_full_140423305666456: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305666456: core_fifo_inputs_t;
        signal outputs_full_140423305666456: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305666512: core_fifo_inputs_t;
        signal fifo_full_140423305666512: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305666512: core_fifo_inputs_t;
        signal outputs_full_140423305666512: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305674824: core_fifo_inputs_t;
        signal fifo_full_140423305674824: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305674824: core_fifo_inputs_t;
        signal outputs_full_140423305674824: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305674880: core_fifo_inputs_t;
        signal fifo_full_140423305674880: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305674880: core_fifo_inputs_t;
        signal outputs_full_140423305674880: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305674936: core_fifo_inputs_t;
        signal fifo_full_140423305674936: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305674936: core_fifo_inputs_t;
        signal outputs_full_140423305674936: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305674992: core_fifo_inputs_t;
        signal fifo_full_140423305674992: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305674992: core_fifo_inputs_t;
        signal outputs_full_140423305674992: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305675048: core_fifo_inputs_t;
        signal fifo_full_140423305675048: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305675048: core_fifo_inputs_t;
        signal outputs_full_140423305675048: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305675104: core_fifo_inputs_t;
        signal fifo_full_140423305675104: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305675104: core_fifo_inputs_t;
        signal outputs_full_140423305675104: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305675160: core_fifo_inputs_t;
        signal fifo_full_140423305675160: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305675160: core_fifo_inputs_t;
        signal outputs_full_140423305675160: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305675216: core_fifo_inputs_t;
        signal fifo_full_140423305675216: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305675216: core_fifo_inputs_t;
        signal outputs_full_140423305675216: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305675272: core_fifo_inputs_t;
        signal fifo_full_140423305675272: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305675272: core_fifo_inputs_t;
        signal outputs_full_140423305675272: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305675328: core_fifo_inputs_t;
        signal fifo_full_140423305675328: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305675328: core_fifo_inputs_t;
        signal outputs_full_140423305675328: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305675384: core_fifo_inputs_t;
        signal fifo_full_140423305675384: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305675384: core_fifo_inputs_t;
        signal outputs_full_140423305675384: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305675440: core_fifo_inputs_t;
        signal fifo_full_140423305675440: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305675440: core_fifo_inputs_t;
        signal outputs_full_140423305675440: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305675496: core_fifo_inputs_t;
        signal fifo_full_140423305675496: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305675496: core_fifo_inputs_t;
        signal outputs_full_140423305675496: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305675552: core_fifo_inputs_t;
        signal fifo_full_140423305675552: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305675552: core_fifo_inputs_t;
        signal outputs_full_140423305675552: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305675608: core_fifo_inputs_t;
        signal fifo_full_140423305675608: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305675608: core_fifo_inputs_t;
        signal outputs_full_140423305675608: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305675664: core_fifo_inputs_t;
        signal fifo_full_140423305675664: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305675664: core_fifo_inputs_t;
        signal outputs_full_140423305675664: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140423305675720: core_fifo_inputs_t;
        signal fifo_full_140423305675720: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140423305675720: core_fifo_inputs_t;
        signal outputs_full_140423305675720: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        

begin
        outputs(0) <= outputs_140423305571464(1);
        outputs_full_140423305571464(1) <= fifo_full(0)

        outputs(1) <= outputs_140423305675720(0);
        outputs_full_140423305675720(0) <= fifo_full(1);
 
    
        fifo_inputs_140423305571408(1) <= outputs_140423305571464(0);
        outputs_full_140423305571464(0) <= fifo_full_140423305571408(1);
        
        fifo_inputs_140423305571632(1) <= outputs_140423305571408(0);
        outputs_full_140423305571408(0) <= fifo_full_140423305571632(1);
        
        fifo_inputs_140423305571464(0) <= outputs_140423305571408(1);
        outputs_full_140423305571408(1) <= fifo_full_140423305571464(0);
        
        fifo_inputs_140423305571688(1) <= outputs_140423305571632(0);
        outputs_full_140423305571632(0) <= fifo_full_140423305571688(1);
        
        fifo_inputs_140423305571408(0) <= outputs_140423305571632(1);
        outputs_full_140423305571632(1) <= fifo_full_140423305571408(0);
        
        fifo_inputs_140423305571744(1) <= outputs_140423305571688(0);
        outputs_full_140423305571688(0) <= fifo_full_140423305571744(1);
        
        fifo_inputs_140423305571632(0) <= outputs_140423305571688(1);
        outputs_full_140423305571688(1) <= fifo_full_140423305571632(0);
        
        fifo_inputs_140423305571576(1) <= outputs_140423305571744(0);
        outputs_full_140423305571744(0) <= fifo_full_140423305571576(1);
        
        fifo_inputs_140423305571688(0) <= outputs_140423305571744(1);
        outputs_full_140423305571744(1) <= fifo_full_140423305571688(0);
        
        fifo_inputs_140423305571800(1) <= outputs_140423305571576(0);
        outputs_full_140423305571576(0) <= fifo_full_140423305571800(1);
        
        fifo_inputs_140423305571744(0) <= outputs_140423305571576(1);
        outputs_full_140423305571576(1) <= fifo_full_140423305571744(0);
        
        fifo_inputs_140423305571856(1) <= outputs_140423305571800(0);
        outputs_full_140423305571800(0) <= fifo_full_140423305571856(1);
        
        fifo_inputs_140423305571576(0) <= outputs_140423305571800(1);
        outputs_full_140423305571800(1) <= fifo_full_140423305571576(0);
        
        fifo_inputs_140423305571912(1) <= outputs_140423305571856(0);
        outputs_full_140423305571856(0) <= fifo_full_140423305571912(1);
        
        fifo_inputs_140423305571800(0) <= outputs_140423305571856(1);
        outputs_full_140423305571856(1) <= fifo_full_140423305571800(0);
        
        fifo_inputs_140423305571968(1) <= outputs_140423305571912(0);
        outputs_full_140423305571912(0) <= fifo_full_140423305571968(1);
        
        fifo_inputs_140423305571856(0) <= outputs_140423305571912(1);
        outputs_full_140423305571912(1) <= fifo_full_140423305571856(0);
        
        fifo_inputs_140423305571520(1) <= outputs_140423305571968(0);
        outputs_full_140423305571968(0) <= fifo_full_140423305571520(1);
        
        fifo_inputs_140423305571912(0) <= outputs_140423305571968(1);
        outputs_full_140423305571968(1) <= fifo_full_140423305571912(0);
        
        fifo_inputs_140423305572024(1) <= outputs_140423305571520(0);
        outputs_full_140423305571520(0) <= fifo_full_140423305572024(1);
        
        fifo_inputs_140423305571968(0) <= outputs_140423305571520(1);
        outputs_full_140423305571520(1) <= fifo_full_140423305571968(0);
        
        fifo_inputs_140423305572080(1) <= outputs_140423305572024(0);
        outputs_full_140423305572024(0) <= fifo_full_140423305572080(1);
        
        fifo_inputs_140423305571520(0) <= outputs_140423305572024(1);
        outputs_full_140423305572024(1) <= fifo_full_140423305571520(0);
        
        fifo_inputs_140423305572136(1) <= outputs_140423305572080(0);
        outputs_full_140423305572080(0) <= fifo_full_140423305572136(1);
        
        fifo_inputs_140423305572024(0) <= outputs_140423305572080(1);
        outputs_full_140423305572080(1) <= fifo_full_140423305572024(0);
        
        fifo_inputs_140423305572192(1) <= outputs_140423305572136(0);
        outputs_full_140423305572136(0) <= fifo_full_140423305572192(1);
        
        fifo_inputs_140423305572080(0) <= outputs_140423305572136(1);
        outputs_full_140423305572136(1) <= fifo_full_140423305572080(0);
        
        fifo_inputs_140423305572248(1) <= outputs_140423305572192(0);
        outputs_full_140423305572192(0) <= fifo_full_140423305572248(1);
        
        fifo_inputs_140423305572136(0) <= outputs_140423305572192(1);
        outputs_full_140423305572192(1) <= fifo_full_140423305572136(0);
        
        fifo_inputs_140423305572304(1) <= outputs_140423305572248(0);
        outputs_full_140423305572248(0) <= fifo_full_140423305572304(1);
        
        fifo_inputs_140423305572192(0) <= outputs_140423305572248(1);
        outputs_full_140423305572248(1) <= fifo_full_140423305572192(0);
        
        fifo_inputs_140423305621576(1) <= outputs_140423305572304(0);
        outputs_full_140423305572304(0) <= fifo_full_140423305621576(1);
        
        fifo_inputs_140423305572248(0) <= outputs_140423305572304(1);
        outputs_full_140423305572304(1) <= fifo_full_140423305572248(0);
        
        fifo_inputs_140423305621632(1) <= outputs_140423305621576(0);
        outputs_full_140423305621576(0) <= fifo_full_140423305621632(1);
        
        fifo_inputs_140423305572304(0) <= outputs_140423305621576(1);
        outputs_full_140423305621576(1) <= fifo_full_140423305572304(0);
        
        fifo_inputs_140423305621688(1) <= outputs_140423305621632(0);
        outputs_full_140423305621632(0) <= fifo_full_140423305621688(1);
        
        fifo_inputs_140423305621576(0) <= outputs_140423305621632(1);
        outputs_full_140423305621632(1) <= fifo_full_140423305621576(0);
        
        fifo_inputs_140423305621744(1) <= outputs_140423305621688(0);
        outputs_full_140423305621688(0) <= fifo_full_140423305621744(1);
        
        fifo_inputs_140423305621632(0) <= outputs_140423305621688(1);
        outputs_full_140423305621688(1) <= fifo_full_140423305621632(0);
        
        fifo_inputs_140423305621800(1) <= outputs_140423305621744(0);
        outputs_full_140423305621744(0) <= fifo_full_140423305621800(1);
        
        fifo_inputs_140423305621688(0) <= outputs_140423305621744(1);
        outputs_full_140423305621744(1) <= fifo_full_140423305621688(0);
        
        fifo_inputs_140423305621856(1) <= outputs_140423305621800(0);
        outputs_full_140423305621800(0) <= fifo_full_140423305621856(1);
        
        fifo_inputs_140423305621744(0) <= outputs_140423305621800(1);
        outputs_full_140423305621800(1) <= fifo_full_140423305621744(0);
        
        fifo_inputs_140423305621912(1) <= outputs_140423305621856(0);
        outputs_full_140423305621856(0) <= fifo_full_140423305621912(1);
        
        fifo_inputs_140423305621800(0) <= outputs_140423305621856(1);
        outputs_full_140423305621856(1) <= fifo_full_140423305621800(0);
        
        fifo_inputs_140423305621968(1) <= outputs_140423305621912(0);
        outputs_full_140423305621912(0) <= fifo_full_140423305621968(1);
        
        fifo_inputs_140423305621856(0) <= outputs_140423305621912(1);
        outputs_full_140423305621912(1) <= fifo_full_140423305621856(0);
        
        fifo_inputs_140423305622024(1) <= outputs_140423305621968(0);
        outputs_full_140423305621968(0) <= fifo_full_140423305622024(1);
        
        fifo_inputs_140423305621912(0) <= outputs_140423305621968(1);
        outputs_full_140423305621968(1) <= fifo_full_140423305621912(0);
        
        fifo_inputs_140423305622080(1) <= outputs_140423305622024(0);
        outputs_full_140423305622024(0) <= fifo_full_140423305622080(1);
        
        fifo_inputs_140423305621968(0) <= outputs_140423305622024(1);
        outputs_full_140423305622024(1) <= fifo_full_140423305621968(0);
        
        fifo_inputs_140423305622136(1) <= outputs_140423305622080(0);
        outputs_full_140423305622080(0) <= fifo_full_140423305622136(1);
        
        fifo_inputs_140423305622024(0) <= outputs_140423305622080(1);
        outputs_full_140423305622080(1) <= fifo_full_140423305622024(0);
        
        fifo_inputs_140423305622192(1) <= outputs_140423305622136(0);
        outputs_full_140423305622136(0) <= fifo_full_140423305622192(1);
        
        fifo_inputs_140423305622080(0) <= outputs_140423305622136(1);
        outputs_full_140423305622136(1) <= fifo_full_140423305622080(0);
        
        fifo_inputs_140423305622248(1) <= outputs_140423305622192(0);
        outputs_full_140423305622192(0) <= fifo_full_140423305622248(1);
        
        fifo_inputs_140423305622136(0) <= outputs_140423305622192(1);
        outputs_full_140423305622192(1) <= fifo_full_140423305622136(0);
        
        fifo_inputs_140423305622304(1) <= outputs_140423305622248(0);
        outputs_full_140423305622248(0) <= fifo_full_140423305622304(1);
        
        fifo_inputs_140423305622192(0) <= outputs_140423305622248(1);
        outputs_full_140423305622248(1) <= fifo_full_140423305622192(0);
        
        fifo_inputs_140423305622360(1) <= outputs_140423305622304(0);
        outputs_full_140423305622304(0) <= fifo_full_140423305622360(1);
        
        fifo_inputs_140423305622248(0) <= outputs_140423305622304(1);
        outputs_full_140423305622304(1) <= fifo_full_140423305622248(0);
        
        fifo_inputs_140423305622416(1) <= outputs_140423305622360(0);
        outputs_full_140423305622360(0) <= fifo_full_140423305622416(1);
        
        fifo_inputs_140423305622304(0) <= outputs_140423305622360(1);
        outputs_full_140423305622360(1) <= fifo_full_140423305622304(0);
        
        fifo_inputs_140423305622472(1) <= outputs_140423305622416(0);
        outputs_full_140423305622416(0) <= fifo_full_140423305622472(1);
        
        fifo_inputs_140423305622360(0) <= outputs_140423305622416(1);
        outputs_full_140423305622416(1) <= fifo_full_140423305622360(0);
        
        fifo_inputs_140423305622528(1) <= outputs_140423305622472(0);
        outputs_full_140423305622472(0) <= fifo_full_140423305622528(1);
        
        fifo_inputs_140423305622416(0) <= outputs_140423305622472(1);
        outputs_full_140423305622472(1) <= fifo_full_140423305622416(0);
        
        fifo_inputs_140423305622584(1) <= outputs_140423305622528(0);
        outputs_full_140423305622528(0) <= fifo_full_140423305622584(1);
        
        fifo_inputs_140423305622472(0) <= outputs_140423305622528(1);
        outputs_full_140423305622528(1) <= fifo_full_140423305622472(0);
        
        fifo_inputs_140423305622640(1) <= outputs_140423305622584(0);
        outputs_full_140423305622584(0) <= fifo_full_140423305622640(1);
        
        fifo_inputs_140423305622528(0) <= outputs_140423305622584(1);
        outputs_full_140423305622584(1) <= fifo_full_140423305622528(0);
        
        fifo_inputs_140423305622696(1) <= outputs_140423305622640(0);
        outputs_full_140423305622640(0) <= fifo_full_140423305622696(1);
        
        fifo_inputs_140423305622584(0) <= outputs_140423305622640(1);
        outputs_full_140423305622640(1) <= fifo_full_140423305622584(0);
        
        fifo_inputs_140423305622752(1) <= outputs_140423305622696(0);
        outputs_full_140423305622696(0) <= fifo_full_140423305622752(1);
        
        fifo_inputs_140423305622640(0) <= outputs_140423305622696(1);
        outputs_full_140423305622696(1) <= fifo_full_140423305622640(0);
        
        fifo_inputs_140423305622808(1) <= outputs_140423305622752(0);
        outputs_full_140423305622752(0) <= fifo_full_140423305622808(1);
        
        fifo_inputs_140423305622696(0) <= outputs_140423305622752(1);
        outputs_full_140423305622752(1) <= fifo_full_140423305622696(0);
        
        fifo_inputs_140423305622864(1) <= outputs_140423305622808(0);
        outputs_full_140423305622808(0) <= fifo_full_140423305622864(1);
        
        fifo_inputs_140423305622752(0) <= outputs_140423305622808(1);
        outputs_full_140423305622808(1) <= fifo_full_140423305622752(0);
        
        fifo_inputs_140423305622920(1) <= outputs_140423305622864(0);
        outputs_full_140423305622864(0) <= fifo_full_140423305622920(1);
        
        fifo_inputs_140423305622808(0) <= outputs_140423305622864(1);
        outputs_full_140423305622864(1) <= fifo_full_140423305622808(0);
        
        fifo_inputs_140423305622976(1) <= outputs_140423305622920(0);
        outputs_full_140423305622920(0) <= fifo_full_140423305622976(1);
        
        fifo_inputs_140423305622864(0) <= outputs_140423305622920(1);
        outputs_full_140423305622920(1) <= fifo_full_140423305622864(0);
        
        fifo_inputs_140423305623032(1) <= outputs_140423305622976(0);
        outputs_full_140423305622976(0) <= fifo_full_140423305623032(1);
        
        fifo_inputs_140423305622920(0) <= outputs_140423305622976(1);
        outputs_full_140423305622976(1) <= fifo_full_140423305622920(0);
        
        fifo_inputs_140423305623088(1) <= outputs_140423305623032(0);
        outputs_full_140423305623032(0) <= fifo_full_140423305623088(1);
        
        fifo_inputs_140423305622976(0) <= outputs_140423305623032(1);
        outputs_full_140423305623032(1) <= fifo_full_140423305622976(0);
        
        fifo_inputs_140423305623144(1) <= outputs_140423305623088(0);
        outputs_full_140423305623088(0) <= fifo_full_140423305623144(1);
        
        fifo_inputs_140423305623032(0) <= outputs_140423305623088(1);
        outputs_full_140423305623088(1) <= fifo_full_140423305623032(0);
        
        fifo_inputs_140423305623200(1) <= outputs_140423305623144(0);
        outputs_full_140423305623144(0) <= fifo_full_140423305623200(1);
        
        fifo_inputs_140423305623088(0) <= outputs_140423305623144(1);
        outputs_full_140423305623144(1) <= fifo_full_140423305623088(0);
        
        fifo_inputs_140423305623256(1) <= outputs_140423305623200(0);
        outputs_full_140423305623200(0) <= fifo_full_140423305623256(1);
        
        fifo_inputs_140423305623144(0) <= outputs_140423305623200(1);
        outputs_full_140423305623200(1) <= fifo_full_140423305623144(0);
        
        fifo_inputs_140423305623312(1) <= outputs_140423305623256(0);
        outputs_full_140423305623256(0) <= fifo_full_140423305623312(1);
        
        fifo_inputs_140423305623200(0) <= outputs_140423305623256(1);
        outputs_full_140423305623256(1) <= fifo_full_140423305623200(0);
        
        fifo_inputs_140423305623368(1) <= outputs_140423305623312(0);
        outputs_full_140423305623312(0) <= fifo_full_140423305623368(1);
        
        fifo_inputs_140423305623256(0) <= outputs_140423305623312(1);
        outputs_full_140423305623312(1) <= fifo_full_140423305623256(0);
        
        fifo_inputs_140423305623424(1) <= outputs_140423305623368(0);
        outputs_full_140423305623368(0) <= fifo_full_140423305623424(1);
        
        fifo_inputs_140423305623312(0) <= outputs_140423305623368(1);
        outputs_full_140423305623368(1) <= fifo_full_140423305623312(0);
        
        fifo_inputs_140423305623480(1) <= outputs_140423305623424(0);
        outputs_full_140423305623424(0) <= fifo_full_140423305623480(1);
        
        fifo_inputs_140423305623368(0) <= outputs_140423305623424(1);
        outputs_full_140423305623424(1) <= fifo_full_140423305623368(0);
        
        fifo_inputs_140423305623536(1) <= outputs_140423305623480(0);
        outputs_full_140423305623480(0) <= fifo_full_140423305623536(1);
        
        fifo_inputs_140423305623424(0) <= outputs_140423305623480(1);
        outputs_full_140423305623480(1) <= fifo_full_140423305623424(0);
        
        fifo_inputs_140423305623592(1) <= outputs_140423305623536(0);
        outputs_full_140423305623536(0) <= fifo_full_140423305623592(1);
        
        fifo_inputs_140423305623480(0) <= outputs_140423305623536(1);
        outputs_full_140423305623536(1) <= fifo_full_140423305623480(0);
        
        fifo_inputs_140423305623648(1) <= outputs_140423305623592(0);
        outputs_full_140423305623592(0) <= fifo_full_140423305623648(1);
        
        fifo_inputs_140423305623536(0) <= outputs_140423305623592(1);
        outputs_full_140423305623592(1) <= fifo_full_140423305623536(0);
        
        fifo_inputs_140423305623704(1) <= outputs_140423305623648(0);
        outputs_full_140423305623648(0) <= fifo_full_140423305623704(1);
        
        fifo_inputs_140423305623592(0) <= outputs_140423305623648(1);
        outputs_full_140423305623648(1) <= fifo_full_140423305623592(0);
        
        fifo_inputs_140423305623760(1) <= outputs_140423305623704(0);
        outputs_full_140423305623704(0) <= fifo_full_140423305623760(1);
        
        fifo_inputs_140423305623648(0) <= outputs_140423305623704(1);
        outputs_full_140423305623704(1) <= fifo_full_140423305623648(0);
        
        fifo_inputs_140423305623816(1) <= outputs_140423305623760(0);
        outputs_full_140423305623760(0) <= fifo_full_140423305623816(1);
        
        fifo_inputs_140423305623704(0) <= outputs_140423305623760(1);
        outputs_full_140423305623760(1) <= fifo_full_140423305623704(0);
        
        fifo_inputs_140423305623872(1) <= outputs_140423305623816(0);
        outputs_full_140423305623816(0) <= fifo_full_140423305623872(1);
        
        fifo_inputs_140423305623760(0) <= outputs_140423305623816(1);
        outputs_full_140423305623816(1) <= fifo_full_140423305623760(0);
        
        fifo_inputs_140423305623928(1) <= outputs_140423305623872(0);
        outputs_full_140423305623872(0) <= fifo_full_140423305623928(1);
        
        fifo_inputs_140423305623816(0) <= outputs_140423305623872(1);
        outputs_full_140423305623872(1) <= fifo_full_140423305623816(0);
        
        fifo_inputs_140423305623984(1) <= outputs_140423305623928(0);
        outputs_full_140423305623928(0) <= fifo_full_140423305623984(1);
        
        fifo_inputs_140423305623872(0) <= outputs_140423305623928(1);
        outputs_full_140423305623928(1) <= fifo_full_140423305623872(0);
        
        fifo_inputs_140423305624040(1) <= outputs_140423305623984(0);
        outputs_full_140423305623984(0) <= fifo_full_140423305624040(1);
        
        fifo_inputs_140423305623928(0) <= outputs_140423305623984(1);
        outputs_full_140423305623984(1) <= fifo_full_140423305623928(0);
        
        fifo_inputs_140423305624096(1) <= outputs_140423305624040(0);
        outputs_full_140423305624040(0) <= fifo_full_140423305624096(1);
        
        fifo_inputs_140423305623984(0) <= outputs_140423305624040(1);
        outputs_full_140423305624040(1) <= fifo_full_140423305623984(0);
        
        fifo_inputs_140423305624152(1) <= outputs_140423305624096(0);
        outputs_full_140423305624096(0) <= fifo_full_140423305624152(1);
        
        fifo_inputs_140423305624040(0) <= outputs_140423305624096(1);
        outputs_full_140423305624096(1) <= fifo_full_140423305624040(0);
        
        fifo_inputs_140423305624208(1) <= outputs_140423305624152(0);
        outputs_full_140423305624152(0) <= fifo_full_140423305624208(1);
        
        fifo_inputs_140423305624096(0) <= outputs_140423305624152(1);
        outputs_full_140423305624152(1) <= fifo_full_140423305624096(0);
        
        fifo_inputs_140423305624264(1) <= outputs_140423305624208(0);
        outputs_full_140423305624208(0) <= fifo_full_140423305624264(1);
        
        fifo_inputs_140423305624152(0) <= outputs_140423305624208(1);
        outputs_full_140423305624208(1) <= fifo_full_140423305624152(0);
        
        fifo_inputs_140423305624320(1) <= outputs_140423305624264(0);
        outputs_full_140423305624264(0) <= fifo_full_140423305624320(1);
        
        fifo_inputs_140423305624208(0) <= outputs_140423305624264(1);
        outputs_full_140423305624264(1) <= fifo_full_140423305624208(0);
        
        fifo_inputs_140423305624376(1) <= outputs_140423305624320(0);
        outputs_full_140423305624320(0) <= fifo_full_140423305624376(1);
        
        fifo_inputs_140423305624264(0) <= outputs_140423305624320(1);
        outputs_full_140423305624320(1) <= fifo_full_140423305624264(0);
        
        fifo_inputs_140423305624432(1) <= outputs_140423305624376(0);
        outputs_full_140423305624376(0) <= fifo_full_140423305624432(1);
        
        fifo_inputs_140423305624320(0) <= outputs_140423305624376(1);
        outputs_full_140423305624376(1) <= fifo_full_140423305624320(0);
        
        fifo_inputs_140423305624488(1) <= outputs_140423305624432(0);
        outputs_full_140423305624432(0) <= fifo_full_140423305624488(1);
        
        fifo_inputs_140423305624376(0) <= outputs_140423305624432(1);
        outputs_full_140423305624432(1) <= fifo_full_140423305624376(0);
        
        fifo_inputs_140423305624544(1) <= outputs_140423305624488(0);
        outputs_full_140423305624488(0) <= fifo_full_140423305624544(1);
        
        fifo_inputs_140423305624432(0) <= outputs_140423305624488(1);
        outputs_full_140423305624488(1) <= fifo_full_140423305624432(0);
        
        fifo_inputs_140423305624600(1) <= outputs_140423305624544(0);
        outputs_full_140423305624544(0) <= fifo_full_140423305624600(1);
        
        fifo_inputs_140423305624488(0) <= outputs_140423305624544(1);
        outputs_full_140423305624544(1) <= fifo_full_140423305624488(0);
        
        fifo_inputs_140423305624656(1) <= outputs_140423305624600(0);
        outputs_full_140423305624600(0) <= fifo_full_140423305624656(1);
        
        fifo_inputs_140423305624544(0) <= outputs_140423305624600(1);
        outputs_full_140423305624600(1) <= fifo_full_140423305624544(0);
        
        fifo_inputs_140423305624712(1) <= outputs_140423305624656(0);
        outputs_full_140423305624656(0) <= fifo_full_140423305624712(1);
        
        fifo_inputs_140423305624600(0) <= outputs_140423305624656(1);
        outputs_full_140423305624656(1) <= fifo_full_140423305624600(0);
        
        fifo_inputs_140423305624768(1) <= outputs_140423305624712(0);
        outputs_full_140423305624712(0) <= fifo_full_140423305624768(1);
        
        fifo_inputs_140423305624656(0) <= outputs_140423305624712(1);
        outputs_full_140423305624712(1) <= fifo_full_140423305624656(0);
        
        fifo_inputs_140423305624824(1) <= outputs_140423305624768(0);
        outputs_full_140423305624768(0) <= fifo_full_140423305624824(1);
        
        fifo_inputs_140423305624712(0) <= outputs_140423305624768(1);
        outputs_full_140423305624768(1) <= fifo_full_140423305624712(0);
        
        fifo_inputs_140423305624880(1) <= outputs_140423305624824(0);
        outputs_full_140423305624824(0) <= fifo_full_140423305624880(1);
        
        fifo_inputs_140423305624768(0) <= outputs_140423305624824(1);
        outputs_full_140423305624824(1) <= fifo_full_140423305624768(0);
        
        fifo_inputs_140423305624936(1) <= outputs_140423305624880(0);
        outputs_full_140423305624880(0) <= fifo_full_140423305624936(1);
        
        fifo_inputs_140423305624824(0) <= outputs_140423305624880(1);
        outputs_full_140423305624880(1) <= fifo_full_140423305624824(0);
        
        fifo_inputs_140423305624992(1) <= outputs_140423305624936(0);
        outputs_full_140423305624936(0) <= fifo_full_140423305624992(1);
        
        fifo_inputs_140423305624880(0) <= outputs_140423305624936(1);
        outputs_full_140423305624936(1) <= fifo_full_140423305624880(0);
        
        fifo_inputs_140423305625048(1) <= outputs_140423305624992(0);
        outputs_full_140423305624992(0) <= fifo_full_140423305625048(1);
        
        fifo_inputs_140423305624936(0) <= outputs_140423305624992(1);
        outputs_full_140423305624992(1) <= fifo_full_140423305624936(0);
        
        fifo_inputs_140423305625104(1) <= outputs_140423305625048(0);
        outputs_full_140423305625048(0) <= fifo_full_140423305625104(1);
        
        fifo_inputs_140423305624992(0) <= outputs_140423305625048(1);
        outputs_full_140423305625048(1) <= fifo_full_140423305624992(0);
        
        fifo_inputs_140423305625160(1) <= outputs_140423305625104(0);
        outputs_full_140423305625104(0) <= fifo_full_140423305625160(1);
        
        fifo_inputs_140423305625048(0) <= outputs_140423305625104(1);
        outputs_full_140423305625104(1) <= fifo_full_140423305625048(0);
        
        fifo_inputs_140423305625216(1) <= outputs_140423305625160(0);
        outputs_full_140423305625160(0) <= fifo_full_140423305625216(1);
        
        fifo_inputs_140423305625104(0) <= outputs_140423305625160(1);
        outputs_full_140423305625160(1) <= fifo_full_140423305625104(0);
        
        fifo_inputs_140423305625272(1) <= outputs_140423305625216(0);
        outputs_full_140423305625216(0) <= fifo_full_140423305625272(1);
        
        fifo_inputs_140423305625160(0) <= outputs_140423305625216(1);
        outputs_full_140423305625216(1) <= fifo_full_140423305625160(0);
        
        fifo_inputs_140423305625328(1) <= outputs_140423305625272(0);
        outputs_full_140423305625272(0) <= fifo_full_140423305625328(1);
        
        fifo_inputs_140423305625216(0) <= outputs_140423305625272(1);
        outputs_full_140423305625272(1) <= fifo_full_140423305625216(0);
        
        fifo_inputs_140423305625384(1) <= outputs_140423305625328(0);
        outputs_full_140423305625328(0) <= fifo_full_140423305625384(1);
        
        fifo_inputs_140423305625272(0) <= outputs_140423305625328(1);
        outputs_full_140423305625328(1) <= fifo_full_140423305625272(0);
        
        fifo_inputs_140423305625440(1) <= outputs_140423305625384(0);
        outputs_full_140423305625384(0) <= fifo_full_140423305625440(1);
        
        fifo_inputs_140423305625328(0) <= outputs_140423305625384(1);
        outputs_full_140423305625384(1) <= fifo_full_140423305625328(0);
        
        fifo_inputs_140423305625496(1) <= outputs_140423305625440(0);
        outputs_full_140423305625440(0) <= fifo_full_140423305625496(1);
        
        fifo_inputs_140423305625384(0) <= outputs_140423305625440(1);
        outputs_full_140423305625440(1) <= fifo_full_140423305625384(0);
        
        fifo_inputs_140423305625552(1) <= outputs_140423305625496(0);
        outputs_full_140423305625496(0) <= fifo_full_140423305625552(1);
        
        fifo_inputs_140423305625440(0) <= outputs_140423305625496(1);
        outputs_full_140423305625496(1) <= fifo_full_140423305625440(0);
        
        fifo_inputs_140423305642056(1) <= outputs_140423305625552(0);
        outputs_full_140423305625552(0) <= fifo_full_140423305642056(1);
        
        fifo_inputs_140423305625496(0) <= outputs_140423305625552(1);
        outputs_full_140423305625552(1) <= fifo_full_140423305625496(0);
        
        fifo_inputs_140423305642112(1) <= outputs_140423305642056(0);
        outputs_full_140423305642056(0) <= fifo_full_140423305642112(1);
        
        fifo_inputs_140423305625552(0) <= outputs_140423305642056(1);
        outputs_full_140423305642056(1) <= fifo_full_140423305625552(0);
        
        fifo_inputs_140423305642168(1) <= outputs_140423305642112(0);
        outputs_full_140423305642112(0) <= fifo_full_140423305642168(1);
        
        fifo_inputs_140423305642056(0) <= outputs_140423305642112(1);
        outputs_full_140423305642112(1) <= fifo_full_140423305642056(0);
        
        fifo_inputs_140423305642224(1) <= outputs_140423305642168(0);
        outputs_full_140423305642168(0) <= fifo_full_140423305642224(1);
        
        fifo_inputs_140423305642112(0) <= outputs_140423305642168(1);
        outputs_full_140423305642168(1) <= fifo_full_140423305642112(0);
        
        fifo_inputs_140423305642280(1) <= outputs_140423305642224(0);
        outputs_full_140423305642224(0) <= fifo_full_140423305642280(1);
        
        fifo_inputs_140423305642168(0) <= outputs_140423305642224(1);
        outputs_full_140423305642224(1) <= fifo_full_140423305642168(0);
        
        fifo_inputs_140423305642336(1) <= outputs_140423305642280(0);
        outputs_full_140423305642280(0) <= fifo_full_140423305642336(1);
        
        fifo_inputs_140423305642224(0) <= outputs_140423305642280(1);
        outputs_full_140423305642280(1) <= fifo_full_140423305642224(0);
        
        fifo_inputs_140423305642392(1) <= outputs_140423305642336(0);
        outputs_full_140423305642336(0) <= fifo_full_140423305642392(1);
        
        fifo_inputs_140423305642280(0) <= outputs_140423305642336(1);
        outputs_full_140423305642336(1) <= fifo_full_140423305642280(0);
        
        fifo_inputs_140423305642448(1) <= outputs_140423305642392(0);
        outputs_full_140423305642392(0) <= fifo_full_140423305642448(1);
        
        fifo_inputs_140423305642336(0) <= outputs_140423305642392(1);
        outputs_full_140423305642392(1) <= fifo_full_140423305642336(0);
        
        fifo_inputs_140423305642504(1) <= outputs_140423305642448(0);
        outputs_full_140423305642448(0) <= fifo_full_140423305642504(1);
        
        fifo_inputs_140423305642392(0) <= outputs_140423305642448(1);
        outputs_full_140423305642448(1) <= fifo_full_140423305642392(0);
        
        fifo_inputs_140423305642560(1) <= outputs_140423305642504(0);
        outputs_full_140423305642504(0) <= fifo_full_140423305642560(1);
        
        fifo_inputs_140423305642448(0) <= outputs_140423305642504(1);
        outputs_full_140423305642504(1) <= fifo_full_140423305642448(0);
        
        fifo_inputs_140423305642616(1) <= outputs_140423305642560(0);
        outputs_full_140423305642560(0) <= fifo_full_140423305642616(1);
        
        fifo_inputs_140423305642504(0) <= outputs_140423305642560(1);
        outputs_full_140423305642560(1) <= fifo_full_140423305642504(0);
        
        fifo_inputs_140423305642672(1) <= outputs_140423305642616(0);
        outputs_full_140423305642616(0) <= fifo_full_140423305642672(1);
        
        fifo_inputs_140423305642560(0) <= outputs_140423305642616(1);
        outputs_full_140423305642616(1) <= fifo_full_140423305642560(0);
        
        fifo_inputs_140423305642728(1) <= outputs_140423305642672(0);
        outputs_full_140423305642672(0) <= fifo_full_140423305642728(1);
        
        fifo_inputs_140423305642616(0) <= outputs_140423305642672(1);
        outputs_full_140423305642672(1) <= fifo_full_140423305642616(0);
        
        fifo_inputs_140423305642784(1) <= outputs_140423305642728(0);
        outputs_full_140423305642728(0) <= fifo_full_140423305642784(1);
        
        fifo_inputs_140423305642672(0) <= outputs_140423305642728(1);
        outputs_full_140423305642728(1) <= fifo_full_140423305642672(0);
        
        fifo_inputs_140423305642840(1) <= outputs_140423305642784(0);
        outputs_full_140423305642784(0) <= fifo_full_140423305642840(1);
        
        fifo_inputs_140423305642728(0) <= outputs_140423305642784(1);
        outputs_full_140423305642784(1) <= fifo_full_140423305642728(0);
        
        fifo_inputs_140423305642896(1) <= outputs_140423305642840(0);
        outputs_full_140423305642840(0) <= fifo_full_140423305642896(1);
        
        fifo_inputs_140423305642784(0) <= outputs_140423305642840(1);
        outputs_full_140423305642840(1) <= fifo_full_140423305642784(0);
        
        fifo_inputs_140423305642952(1) <= outputs_140423305642896(0);
        outputs_full_140423305642896(0) <= fifo_full_140423305642952(1);
        
        fifo_inputs_140423305642840(0) <= outputs_140423305642896(1);
        outputs_full_140423305642896(1) <= fifo_full_140423305642840(0);
        
        fifo_inputs_140423305643008(1) <= outputs_140423305642952(0);
        outputs_full_140423305642952(0) <= fifo_full_140423305643008(1);
        
        fifo_inputs_140423305642896(0) <= outputs_140423305642952(1);
        outputs_full_140423305642952(1) <= fifo_full_140423305642896(0);
        
        fifo_inputs_140423305643064(1) <= outputs_140423305643008(0);
        outputs_full_140423305643008(0) <= fifo_full_140423305643064(1);
        
        fifo_inputs_140423305642952(0) <= outputs_140423305643008(1);
        outputs_full_140423305643008(1) <= fifo_full_140423305642952(0);
        
        fifo_inputs_140423305643120(1) <= outputs_140423305643064(0);
        outputs_full_140423305643064(0) <= fifo_full_140423305643120(1);
        
        fifo_inputs_140423305643008(0) <= outputs_140423305643064(1);
        outputs_full_140423305643064(1) <= fifo_full_140423305643008(0);
        
        fifo_inputs_140423305643176(1) <= outputs_140423305643120(0);
        outputs_full_140423305643120(0) <= fifo_full_140423305643176(1);
        
        fifo_inputs_140423305643064(0) <= outputs_140423305643120(1);
        outputs_full_140423305643120(1) <= fifo_full_140423305643064(0);
        
        fifo_inputs_140423305643232(1) <= outputs_140423305643176(0);
        outputs_full_140423305643176(0) <= fifo_full_140423305643232(1);
        
        fifo_inputs_140423305643120(0) <= outputs_140423305643176(1);
        outputs_full_140423305643176(1) <= fifo_full_140423305643120(0);
        
        fifo_inputs_140423305643288(1) <= outputs_140423305643232(0);
        outputs_full_140423305643232(0) <= fifo_full_140423305643288(1);
        
        fifo_inputs_140423305643176(0) <= outputs_140423305643232(1);
        outputs_full_140423305643232(1) <= fifo_full_140423305643176(0);
        
        fifo_inputs_140423305643344(1) <= outputs_140423305643288(0);
        outputs_full_140423305643288(0) <= fifo_full_140423305643344(1);
        
        fifo_inputs_140423305643232(0) <= outputs_140423305643288(1);
        outputs_full_140423305643288(1) <= fifo_full_140423305643232(0);
        
        fifo_inputs_140423305643400(1) <= outputs_140423305643344(0);
        outputs_full_140423305643344(0) <= fifo_full_140423305643400(1);
        
        fifo_inputs_140423305643288(0) <= outputs_140423305643344(1);
        outputs_full_140423305643344(1) <= fifo_full_140423305643288(0);
        
        fifo_inputs_140423305643456(1) <= outputs_140423305643400(0);
        outputs_full_140423305643400(0) <= fifo_full_140423305643456(1);
        
        fifo_inputs_140423305643344(0) <= outputs_140423305643400(1);
        outputs_full_140423305643400(1) <= fifo_full_140423305643344(0);
        
        fifo_inputs_140423305643512(1) <= outputs_140423305643456(0);
        outputs_full_140423305643456(0) <= fifo_full_140423305643512(1);
        
        fifo_inputs_140423305643400(0) <= outputs_140423305643456(1);
        outputs_full_140423305643456(1) <= fifo_full_140423305643400(0);
        
        fifo_inputs_140423305643568(1) <= outputs_140423305643512(0);
        outputs_full_140423305643512(0) <= fifo_full_140423305643568(1);
        
        fifo_inputs_140423305643456(0) <= outputs_140423305643512(1);
        outputs_full_140423305643512(1) <= fifo_full_140423305643456(0);
        
        fifo_inputs_140423305643624(1) <= outputs_140423305643568(0);
        outputs_full_140423305643568(0) <= fifo_full_140423305643624(1);
        
        fifo_inputs_140423305643512(0) <= outputs_140423305643568(1);
        outputs_full_140423305643568(1) <= fifo_full_140423305643512(0);
        
        fifo_inputs_140423305643680(1) <= outputs_140423305643624(0);
        outputs_full_140423305643624(0) <= fifo_full_140423305643680(1);
        
        fifo_inputs_140423305643568(0) <= outputs_140423305643624(1);
        outputs_full_140423305643624(1) <= fifo_full_140423305643568(0);
        
        fifo_inputs_140423305643736(1) <= outputs_140423305643680(0);
        outputs_full_140423305643680(0) <= fifo_full_140423305643736(1);
        
        fifo_inputs_140423305643624(0) <= outputs_140423305643680(1);
        outputs_full_140423305643680(1) <= fifo_full_140423305643624(0);
        
        fifo_inputs_140423305643792(1) <= outputs_140423305643736(0);
        outputs_full_140423305643736(0) <= fifo_full_140423305643792(1);
        
        fifo_inputs_140423305643680(0) <= outputs_140423305643736(1);
        outputs_full_140423305643736(1) <= fifo_full_140423305643680(0);
        
        fifo_inputs_140423305643848(1) <= outputs_140423305643792(0);
        outputs_full_140423305643792(0) <= fifo_full_140423305643848(1);
        
        fifo_inputs_140423305643736(0) <= outputs_140423305643792(1);
        outputs_full_140423305643792(1) <= fifo_full_140423305643736(0);
        
        fifo_inputs_140423305643904(1) <= outputs_140423305643848(0);
        outputs_full_140423305643848(0) <= fifo_full_140423305643904(1);
        
        fifo_inputs_140423305643792(0) <= outputs_140423305643848(1);
        outputs_full_140423305643848(1) <= fifo_full_140423305643792(0);
        
        fifo_inputs_140423305643960(1) <= outputs_140423305643904(0);
        outputs_full_140423305643904(0) <= fifo_full_140423305643960(1);
        
        fifo_inputs_140423305643848(0) <= outputs_140423305643904(1);
        outputs_full_140423305643904(1) <= fifo_full_140423305643848(0);
        
        fifo_inputs_140423305644016(1) <= outputs_140423305643960(0);
        outputs_full_140423305643960(0) <= fifo_full_140423305644016(1);
        
        fifo_inputs_140423305643904(0) <= outputs_140423305643960(1);
        outputs_full_140423305643960(1) <= fifo_full_140423305643904(0);
        
        fifo_inputs_140423305644072(1) <= outputs_140423305644016(0);
        outputs_full_140423305644016(0) <= fifo_full_140423305644072(1);
        
        fifo_inputs_140423305643960(0) <= outputs_140423305644016(1);
        outputs_full_140423305644016(1) <= fifo_full_140423305643960(0);
        
        fifo_inputs_140423305644128(1) <= outputs_140423305644072(0);
        outputs_full_140423305644072(0) <= fifo_full_140423305644128(1);
        
        fifo_inputs_140423305644016(0) <= outputs_140423305644072(1);
        outputs_full_140423305644072(1) <= fifo_full_140423305644016(0);
        
        fifo_inputs_140423305644184(1) <= outputs_140423305644128(0);
        outputs_full_140423305644128(0) <= fifo_full_140423305644184(1);
        
        fifo_inputs_140423305644072(0) <= outputs_140423305644128(1);
        outputs_full_140423305644128(1) <= fifo_full_140423305644072(0);
        
        fifo_inputs_140423305644240(1) <= outputs_140423305644184(0);
        outputs_full_140423305644184(0) <= fifo_full_140423305644240(1);
        
        fifo_inputs_140423305644128(0) <= outputs_140423305644184(1);
        outputs_full_140423305644184(1) <= fifo_full_140423305644128(0);
        
        fifo_inputs_140423305644296(1) <= outputs_140423305644240(0);
        outputs_full_140423305644240(0) <= fifo_full_140423305644296(1);
        
        fifo_inputs_140423305644184(0) <= outputs_140423305644240(1);
        outputs_full_140423305644240(1) <= fifo_full_140423305644184(0);
        
        fifo_inputs_140423305644352(1) <= outputs_140423305644296(0);
        outputs_full_140423305644296(0) <= fifo_full_140423305644352(1);
        
        fifo_inputs_140423305644240(0) <= outputs_140423305644296(1);
        outputs_full_140423305644296(1) <= fifo_full_140423305644240(0);
        
        fifo_inputs_140423305644408(1) <= outputs_140423305644352(0);
        outputs_full_140423305644352(0) <= fifo_full_140423305644408(1);
        
        fifo_inputs_140423305644296(0) <= outputs_140423305644352(1);
        outputs_full_140423305644352(1) <= fifo_full_140423305644296(0);
        
        fifo_inputs_140423305644464(1) <= outputs_140423305644408(0);
        outputs_full_140423305644408(0) <= fifo_full_140423305644464(1);
        
        fifo_inputs_140423305644352(0) <= outputs_140423305644408(1);
        outputs_full_140423305644408(1) <= fifo_full_140423305644352(0);
        
        fifo_inputs_140423305644520(1) <= outputs_140423305644464(0);
        outputs_full_140423305644464(0) <= fifo_full_140423305644520(1);
        
        fifo_inputs_140423305644408(0) <= outputs_140423305644464(1);
        outputs_full_140423305644464(1) <= fifo_full_140423305644408(0);
        
        fifo_inputs_140423305644576(1) <= outputs_140423305644520(0);
        outputs_full_140423305644520(0) <= fifo_full_140423305644576(1);
        
        fifo_inputs_140423305644464(0) <= outputs_140423305644520(1);
        outputs_full_140423305644520(1) <= fifo_full_140423305644464(0);
        
        fifo_inputs_140423305644632(1) <= outputs_140423305644576(0);
        outputs_full_140423305644576(0) <= fifo_full_140423305644632(1);
        
        fifo_inputs_140423305644520(0) <= outputs_140423305644576(1);
        outputs_full_140423305644576(1) <= fifo_full_140423305644520(0);
        
        fifo_inputs_140423305644688(1) <= outputs_140423305644632(0);
        outputs_full_140423305644632(0) <= fifo_full_140423305644688(1);
        
        fifo_inputs_140423305644576(0) <= outputs_140423305644632(1);
        outputs_full_140423305644632(1) <= fifo_full_140423305644576(0);
        
        fifo_inputs_140423305644744(1) <= outputs_140423305644688(0);
        outputs_full_140423305644688(0) <= fifo_full_140423305644744(1);
        
        fifo_inputs_140423305644632(0) <= outputs_140423305644688(1);
        outputs_full_140423305644688(1) <= fifo_full_140423305644632(0);
        
        fifo_inputs_140423305644800(1) <= outputs_140423305644744(0);
        outputs_full_140423305644744(0) <= fifo_full_140423305644800(1);
        
        fifo_inputs_140423305644688(0) <= outputs_140423305644744(1);
        outputs_full_140423305644744(1) <= fifo_full_140423305644688(0);
        
        fifo_inputs_140423305644856(1) <= outputs_140423305644800(0);
        outputs_full_140423305644800(0) <= fifo_full_140423305644856(1);
        
        fifo_inputs_140423305644744(0) <= outputs_140423305644800(1);
        outputs_full_140423305644800(1) <= fifo_full_140423305644744(0);
        
        fifo_inputs_140423305644912(1) <= outputs_140423305644856(0);
        outputs_full_140423305644856(0) <= fifo_full_140423305644912(1);
        
        fifo_inputs_140423305644800(0) <= outputs_140423305644856(1);
        outputs_full_140423305644856(1) <= fifo_full_140423305644800(0);
        
        fifo_inputs_140423305644968(1) <= outputs_140423305644912(0);
        outputs_full_140423305644912(0) <= fifo_full_140423305644968(1);
        
        fifo_inputs_140423305644856(0) <= outputs_140423305644912(1);
        outputs_full_140423305644912(1) <= fifo_full_140423305644856(0);
        
        fifo_inputs_140423305645024(1) <= outputs_140423305644968(0);
        outputs_full_140423305644968(0) <= fifo_full_140423305645024(1);
        
        fifo_inputs_140423305644912(0) <= outputs_140423305644968(1);
        outputs_full_140423305644968(1) <= fifo_full_140423305644912(0);
        
        fifo_inputs_140423305645080(1) <= outputs_140423305645024(0);
        outputs_full_140423305645024(0) <= fifo_full_140423305645080(1);
        
        fifo_inputs_140423305644968(0) <= outputs_140423305645024(1);
        outputs_full_140423305645024(1) <= fifo_full_140423305644968(0);
        
        fifo_inputs_140423305645136(1) <= outputs_140423305645080(0);
        outputs_full_140423305645080(0) <= fifo_full_140423305645136(1);
        
        fifo_inputs_140423305645024(0) <= outputs_140423305645080(1);
        outputs_full_140423305645080(1) <= fifo_full_140423305645024(0);
        
        fifo_inputs_140423305645192(1) <= outputs_140423305645136(0);
        outputs_full_140423305645136(0) <= fifo_full_140423305645192(1);
        
        fifo_inputs_140423305645080(0) <= outputs_140423305645136(1);
        outputs_full_140423305645136(1) <= fifo_full_140423305645080(0);
        
        fifo_inputs_140423305645248(1) <= outputs_140423305645192(0);
        outputs_full_140423305645192(0) <= fifo_full_140423305645248(1);
        
        fifo_inputs_140423305645136(0) <= outputs_140423305645192(1);
        outputs_full_140423305645192(1) <= fifo_full_140423305645136(0);
        
        fifo_inputs_140423305645304(1) <= outputs_140423305645248(0);
        outputs_full_140423305645248(0) <= fifo_full_140423305645304(1);
        
        fifo_inputs_140423305645192(0) <= outputs_140423305645248(1);
        outputs_full_140423305645248(1) <= fifo_full_140423305645192(0);
        
        fifo_inputs_140423305645360(1) <= outputs_140423305645304(0);
        outputs_full_140423305645304(0) <= fifo_full_140423305645360(1);
        
        fifo_inputs_140423305645248(0) <= outputs_140423305645304(1);
        outputs_full_140423305645304(1) <= fifo_full_140423305645248(0);
        
        fifo_inputs_140423305645416(1) <= outputs_140423305645360(0);
        outputs_full_140423305645360(0) <= fifo_full_140423305645416(1);
        
        fifo_inputs_140423305645304(0) <= outputs_140423305645360(1);
        outputs_full_140423305645360(1) <= fifo_full_140423305645304(0);
        
        fifo_inputs_140423305645472(1) <= outputs_140423305645416(0);
        outputs_full_140423305645416(0) <= fifo_full_140423305645472(1);
        
        fifo_inputs_140423305645360(0) <= outputs_140423305645416(1);
        outputs_full_140423305645416(1) <= fifo_full_140423305645360(0);
        
        fifo_inputs_140423305645528(1) <= outputs_140423305645472(0);
        outputs_full_140423305645472(0) <= fifo_full_140423305645528(1);
        
        fifo_inputs_140423305645416(0) <= outputs_140423305645472(1);
        outputs_full_140423305645472(1) <= fifo_full_140423305645416(0);
        
        fifo_inputs_140423305645584(1) <= outputs_140423305645528(0);
        outputs_full_140423305645528(0) <= fifo_full_140423305645584(1);
        
        fifo_inputs_140423305645472(0) <= outputs_140423305645528(1);
        outputs_full_140423305645528(1) <= fifo_full_140423305645472(0);
        
        fifo_inputs_140423305645640(1) <= outputs_140423305645584(0);
        outputs_full_140423305645584(0) <= fifo_full_140423305645640(1);
        
        fifo_inputs_140423305645528(0) <= outputs_140423305645584(1);
        outputs_full_140423305645584(1) <= fifo_full_140423305645528(0);
        
        fifo_inputs_140423329706112(1) <= outputs_140423305645640(0);
        outputs_full_140423305645640(0) <= fifo_full_140423329706112(1);
        
        fifo_inputs_140423305645584(0) <= outputs_140423305645640(1);
        outputs_full_140423305645640(1) <= fifo_full_140423305645584(0);
        
        fifo_inputs_140423305571240(1) <= outputs_140423329706112(0);
        outputs_full_140423329706112(0) <= fifo_full_140423305571240(1);
        
        fifo_inputs_140423305645640(0) <= outputs_140423329706112(1);
        outputs_full_140423329706112(1) <= fifo_full_140423305645640(0);
        
        fifo_inputs_140423305571016(1) <= outputs_140423305571240(0);
        outputs_full_140423305571240(0) <= fifo_full_140423305571016(1);
        
        fifo_inputs_140423329706112(0) <= outputs_140423305571240(1);
        outputs_full_140423305571240(1) <= fifo_full_140423329706112(0);
        
        fifo_inputs_140423305571296(1) <= outputs_140423305571016(0);
        outputs_full_140423305571016(0) <= fifo_full_140423305571296(1);
        
        fifo_inputs_140423305571240(0) <= outputs_140423305571016(1);
        outputs_full_140423305571016(1) <= fifo_full_140423305571240(0);
        
        fifo_inputs_140423305571072(1) <= outputs_140423305571296(0);
        outputs_full_140423305571296(0) <= fifo_full_140423305571072(1);
        
        fifo_inputs_140423305571016(0) <= outputs_140423305571296(1);
        outputs_full_140423305571296(1) <= fifo_full_140423305571016(0);
        
        fifo_inputs_140423305571128(1) <= outputs_140423305571072(0);
        outputs_full_140423305571072(0) <= fifo_full_140423305571128(1);
        
        fifo_inputs_140423305571296(0) <= outputs_140423305571072(1);
        outputs_full_140423305571072(1) <= fifo_full_140423305571296(0);
        
        fifo_inputs_140423305645696(1) <= outputs_140423305571128(0);
        outputs_full_140423305571128(0) <= fifo_full_140423305645696(1);
        
        fifo_inputs_140423305571072(0) <= outputs_140423305571128(1);
        outputs_full_140423305571128(1) <= fifo_full_140423305571072(0);
        
        fifo_inputs_140423305645752(1) <= outputs_140423305645696(0);
        outputs_full_140423305645696(0) <= fifo_full_140423305645752(1);
        
        fifo_inputs_140423305571128(0) <= outputs_140423305645696(1);
        outputs_full_140423305645696(1) <= fifo_full_140423305571128(0);
        
        fifo_inputs_140423305645808(1) <= outputs_140423305645752(0);
        outputs_full_140423305645752(0) <= fifo_full_140423305645808(1);
        
        fifo_inputs_140423305645696(0) <= outputs_140423305645752(1);
        outputs_full_140423305645752(1) <= fifo_full_140423305645696(0);
        
        fifo_inputs_140423305645864(1) <= outputs_140423305645808(0);
        outputs_full_140423305645808(0) <= fifo_full_140423305645864(1);
        
        fifo_inputs_140423305645752(0) <= outputs_140423305645808(1);
        outputs_full_140423305645808(1) <= fifo_full_140423305645752(0);
        
        fifo_inputs_140423305645920(1) <= outputs_140423305645864(0);
        outputs_full_140423305645864(0) <= fifo_full_140423305645920(1);
        
        fifo_inputs_140423305645808(0) <= outputs_140423305645864(1);
        outputs_full_140423305645864(1) <= fifo_full_140423305645808(0);
        
        fifo_inputs_140423305645976(1) <= outputs_140423305645920(0);
        outputs_full_140423305645920(0) <= fifo_full_140423305645976(1);
        
        fifo_inputs_140423305645864(0) <= outputs_140423305645920(1);
        outputs_full_140423305645920(1) <= fifo_full_140423305645864(0);
        
        fifo_inputs_140423305646032(1) <= outputs_140423305645976(0);
        outputs_full_140423305645976(0) <= fifo_full_140423305646032(1);
        
        fifo_inputs_140423305645920(0) <= outputs_140423305645976(1);
        outputs_full_140423305645976(1) <= fifo_full_140423305645920(0);
        
        fifo_inputs_140423305662536(1) <= outputs_140423305646032(0);
        outputs_full_140423305646032(0) <= fifo_full_140423305662536(1);
        
        fifo_inputs_140423305645976(0) <= outputs_140423305646032(1);
        outputs_full_140423305646032(1) <= fifo_full_140423305645976(0);
        
        fifo_inputs_140423305662592(1) <= outputs_140423305662536(0);
        outputs_full_140423305662536(0) <= fifo_full_140423305662592(1);
        
        fifo_inputs_140423305646032(0) <= outputs_140423305662536(1);
        outputs_full_140423305662536(1) <= fifo_full_140423305646032(0);
        
        fifo_inputs_140423305662648(1) <= outputs_140423305662592(0);
        outputs_full_140423305662592(0) <= fifo_full_140423305662648(1);
        
        fifo_inputs_140423305662536(0) <= outputs_140423305662592(1);
        outputs_full_140423305662592(1) <= fifo_full_140423305662536(0);
        
        fifo_inputs_140423305662704(1) <= outputs_140423305662648(0);
        outputs_full_140423305662648(0) <= fifo_full_140423305662704(1);
        
        fifo_inputs_140423305662592(0) <= outputs_140423305662648(1);
        outputs_full_140423305662648(1) <= fifo_full_140423305662592(0);
        
        fifo_inputs_140423305662760(1) <= outputs_140423305662704(0);
        outputs_full_140423305662704(0) <= fifo_full_140423305662760(1);
        
        fifo_inputs_140423305662648(0) <= outputs_140423305662704(1);
        outputs_full_140423305662704(1) <= fifo_full_140423305662648(0);
        
        fifo_inputs_140423305662816(1) <= outputs_140423305662760(0);
        outputs_full_140423305662760(0) <= fifo_full_140423305662816(1);
        
        fifo_inputs_140423305662704(0) <= outputs_140423305662760(1);
        outputs_full_140423305662760(1) <= fifo_full_140423305662704(0);
        
        fifo_inputs_140423305662872(1) <= outputs_140423305662816(0);
        outputs_full_140423305662816(0) <= fifo_full_140423305662872(1);
        
        fifo_inputs_140423305662760(0) <= outputs_140423305662816(1);
        outputs_full_140423305662816(1) <= fifo_full_140423305662760(0);
        
        fifo_inputs_140423305662928(1) <= outputs_140423305662872(0);
        outputs_full_140423305662872(0) <= fifo_full_140423305662928(1);
        
        fifo_inputs_140423305662816(0) <= outputs_140423305662872(1);
        outputs_full_140423305662872(1) <= fifo_full_140423305662816(0);
        
        fifo_inputs_140423305662984(1) <= outputs_140423305662928(0);
        outputs_full_140423305662928(0) <= fifo_full_140423305662984(1);
        
        fifo_inputs_140423305662872(0) <= outputs_140423305662928(1);
        outputs_full_140423305662928(1) <= fifo_full_140423305662872(0);
        
        fifo_inputs_140423305663040(1) <= outputs_140423305662984(0);
        outputs_full_140423305662984(0) <= fifo_full_140423305663040(1);
        
        fifo_inputs_140423305662928(0) <= outputs_140423305662984(1);
        outputs_full_140423305662984(1) <= fifo_full_140423305662928(0);
        
        fifo_inputs_140423305663096(1) <= outputs_140423305663040(0);
        outputs_full_140423305663040(0) <= fifo_full_140423305663096(1);
        
        fifo_inputs_140423305662984(0) <= outputs_140423305663040(1);
        outputs_full_140423305663040(1) <= fifo_full_140423305662984(0);
        
        fifo_inputs_140423305663152(1) <= outputs_140423305663096(0);
        outputs_full_140423305663096(0) <= fifo_full_140423305663152(1);
        
        fifo_inputs_140423305663040(0) <= outputs_140423305663096(1);
        outputs_full_140423305663096(1) <= fifo_full_140423305663040(0);
        
        fifo_inputs_140423305663208(1) <= outputs_140423305663152(0);
        outputs_full_140423305663152(0) <= fifo_full_140423305663208(1);
        
        fifo_inputs_140423305663096(0) <= outputs_140423305663152(1);
        outputs_full_140423305663152(1) <= fifo_full_140423305663096(0);
        
        fifo_inputs_140423305663264(1) <= outputs_140423305663208(0);
        outputs_full_140423305663208(0) <= fifo_full_140423305663264(1);
        
        fifo_inputs_140423305663152(0) <= outputs_140423305663208(1);
        outputs_full_140423305663208(1) <= fifo_full_140423305663152(0);
        
        fifo_inputs_140423305663320(1) <= outputs_140423305663264(0);
        outputs_full_140423305663264(0) <= fifo_full_140423305663320(1);
        
        fifo_inputs_140423305663208(0) <= outputs_140423305663264(1);
        outputs_full_140423305663264(1) <= fifo_full_140423305663208(0);
        
        fifo_inputs_140423305663376(1) <= outputs_140423305663320(0);
        outputs_full_140423305663320(0) <= fifo_full_140423305663376(1);
        
        fifo_inputs_140423305663264(0) <= outputs_140423305663320(1);
        outputs_full_140423305663320(1) <= fifo_full_140423305663264(0);
        
        fifo_inputs_140423305663432(1) <= outputs_140423305663376(0);
        outputs_full_140423305663376(0) <= fifo_full_140423305663432(1);
        
        fifo_inputs_140423305663320(0) <= outputs_140423305663376(1);
        outputs_full_140423305663376(1) <= fifo_full_140423305663320(0);
        
        fifo_inputs_140423305663488(1) <= outputs_140423305663432(0);
        outputs_full_140423305663432(0) <= fifo_full_140423305663488(1);
        
        fifo_inputs_140423305663376(0) <= outputs_140423305663432(1);
        outputs_full_140423305663432(1) <= fifo_full_140423305663376(0);
        
        fifo_inputs_140423305663544(1) <= outputs_140423305663488(0);
        outputs_full_140423305663488(0) <= fifo_full_140423305663544(1);
        
        fifo_inputs_140423305663432(0) <= outputs_140423305663488(1);
        outputs_full_140423305663488(1) <= fifo_full_140423305663432(0);
        
        fifo_inputs_140423305663600(1) <= outputs_140423305663544(0);
        outputs_full_140423305663544(0) <= fifo_full_140423305663600(1);
        
        fifo_inputs_140423305663488(0) <= outputs_140423305663544(1);
        outputs_full_140423305663544(1) <= fifo_full_140423305663488(0);
        
        fifo_inputs_140423305663656(1) <= outputs_140423305663600(0);
        outputs_full_140423305663600(0) <= fifo_full_140423305663656(1);
        
        fifo_inputs_140423305663544(0) <= outputs_140423305663600(1);
        outputs_full_140423305663600(1) <= fifo_full_140423305663544(0);
        
        fifo_inputs_140423305663712(1) <= outputs_140423305663656(0);
        outputs_full_140423305663656(0) <= fifo_full_140423305663712(1);
        
        fifo_inputs_140423305663600(0) <= outputs_140423305663656(1);
        outputs_full_140423305663656(1) <= fifo_full_140423305663600(0);
        
        fifo_inputs_140423305663768(1) <= outputs_140423305663712(0);
        outputs_full_140423305663712(0) <= fifo_full_140423305663768(1);
        
        fifo_inputs_140423305663656(0) <= outputs_140423305663712(1);
        outputs_full_140423305663712(1) <= fifo_full_140423305663656(0);
        
        fifo_inputs_140423305663824(1) <= outputs_140423305663768(0);
        outputs_full_140423305663768(0) <= fifo_full_140423305663824(1);
        
        fifo_inputs_140423305663712(0) <= outputs_140423305663768(1);
        outputs_full_140423305663768(1) <= fifo_full_140423305663712(0);
        
        fifo_inputs_140423305663880(1) <= outputs_140423305663824(0);
        outputs_full_140423305663824(0) <= fifo_full_140423305663880(1);
        
        fifo_inputs_140423305663768(0) <= outputs_140423305663824(1);
        outputs_full_140423305663824(1) <= fifo_full_140423305663768(0);
        
        fifo_inputs_140423305663936(1) <= outputs_140423305663880(0);
        outputs_full_140423305663880(0) <= fifo_full_140423305663936(1);
        
        fifo_inputs_140423305663824(0) <= outputs_140423305663880(1);
        outputs_full_140423305663880(1) <= fifo_full_140423305663824(0);
        
        fifo_inputs_140423305663992(1) <= outputs_140423305663936(0);
        outputs_full_140423305663936(0) <= fifo_full_140423305663992(1);
        
        fifo_inputs_140423305663880(0) <= outputs_140423305663936(1);
        outputs_full_140423305663936(1) <= fifo_full_140423305663880(0);
        
        fifo_inputs_140423305664048(1) <= outputs_140423305663992(0);
        outputs_full_140423305663992(0) <= fifo_full_140423305664048(1);
        
        fifo_inputs_140423305663936(0) <= outputs_140423305663992(1);
        outputs_full_140423305663992(1) <= fifo_full_140423305663936(0);
        
        fifo_inputs_140423305664104(1) <= outputs_140423305664048(0);
        outputs_full_140423305664048(0) <= fifo_full_140423305664104(1);
        
        fifo_inputs_140423305663992(0) <= outputs_140423305664048(1);
        outputs_full_140423305664048(1) <= fifo_full_140423305663992(0);
        
        fifo_inputs_140423305664160(1) <= outputs_140423305664104(0);
        outputs_full_140423305664104(0) <= fifo_full_140423305664160(1);
        
        fifo_inputs_140423305664048(0) <= outputs_140423305664104(1);
        outputs_full_140423305664104(1) <= fifo_full_140423305664048(0);
        
        fifo_inputs_140423305664216(1) <= outputs_140423305664160(0);
        outputs_full_140423305664160(0) <= fifo_full_140423305664216(1);
        
        fifo_inputs_140423305664104(0) <= outputs_140423305664160(1);
        outputs_full_140423305664160(1) <= fifo_full_140423305664104(0);
        
        fifo_inputs_140423305664272(1) <= outputs_140423305664216(0);
        outputs_full_140423305664216(0) <= fifo_full_140423305664272(1);
        
        fifo_inputs_140423305664160(0) <= outputs_140423305664216(1);
        outputs_full_140423305664216(1) <= fifo_full_140423305664160(0);
        
        fifo_inputs_140423305664328(1) <= outputs_140423305664272(0);
        outputs_full_140423305664272(0) <= fifo_full_140423305664328(1);
        
        fifo_inputs_140423305664216(0) <= outputs_140423305664272(1);
        outputs_full_140423305664272(1) <= fifo_full_140423305664216(0);
        
        fifo_inputs_140423305664384(1) <= outputs_140423305664328(0);
        outputs_full_140423305664328(0) <= fifo_full_140423305664384(1);
        
        fifo_inputs_140423305664272(0) <= outputs_140423305664328(1);
        outputs_full_140423305664328(1) <= fifo_full_140423305664272(0);
        
        fifo_inputs_140423305664440(1) <= outputs_140423305664384(0);
        outputs_full_140423305664384(0) <= fifo_full_140423305664440(1);
        
        fifo_inputs_140423305664328(0) <= outputs_140423305664384(1);
        outputs_full_140423305664384(1) <= fifo_full_140423305664328(0);
        
        fifo_inputs_140423305664496(1) <= outputs_140423305664440(0);
        outputs_full_140423305664440(0) <= fifo_full_140423305664496(1);
        
        fifo_inputs_140423305664384(0) <= outputs_140423305664440(1);
        outputs_full_140423305664440(1) <= fifo_full_140423305664384(0);
        
        fifo_inputs_140423305664552(1) <= outputs_140423305664496(0);
        outputs_full_140423305664496(0) <= fifo_full_140423305664552(1);
        
        fifo_inputs_140423305664440(0) <= outputs_140423305664496(1);
        outputs_full_140423305664496(1) <= fifo_full_140423305664440(0);
        
        fifo_inputs_140423305664608(1) <= outputs_140423305664552(0);
        outputs_full_140423305664552(0) <= fifo_full_140423305664608(1);
        
        fifo_inputs_140423305664496(0) <= outputs_140423305664552(1);
        outputs_full_140423305664552(1) <= fifo_full_140423305664496(0);
        
        fifo_inputs_140423305664664(1) <= outputs_140423305664608(0);
        outputs_full_140423305664608(0) <= fifo_full_140423305664664(1);
        
        fifo_inputs_140423305664552(0) <= outputs_140423305664608(1);
        outputs_full_140423305664608(1) <= fifo_full_140423305664552(0);
        
        fifo_inputs_140423305664720(1) <= outputs_140423305664664(0);
        outputs_full_140423305664664(0) <= fifo_full_140423305664720(1);
        
        fifo_inputs_140423305664608(0) <= outputs_140423305664664(1);
        outputs_full_140423305664664(1) <= fifo_full_140423305664608(0);
        
        fifo_inputs_140423305664776(1) <= outputs_140423305664720(0);
        outputs_full_140423305664720(0) <= fifo_full_140423305664776(1);
        
        fifo_inputs_140423305664664(0) <= outputs_140423305664720(1);
        outputs_full_140423305664720(1) <= fifo_full_140423305664664(0);
        
        fifo_inputs_140423305664832(1) <= outputs_140423305664776(0);
        outputs_full_140423305664776(0) <= fifo_full_140423305664832(1);
        
        fifo_inputs_140423305664720(0) <= outputs_140423305664776(1);
        outputs_full_140423305664776(1) <= fifo_full_140423305664720(0);
        
        fifo_inputs_140423305664888(1) <= outputs_140423305664832(0);
        outputs_full_140423305664832(0) <= fifo_full_140423305664888(1);
        
        fifo_inputs_140423305664776(0) <= outputs_140423305664832(1);
        outputs_full_140423305664832(1) <= fifo_full_140423305664776(0);
        
        fifo_inputs_140423305664944(1) <= outputs_140423305664888(0);
        outputs_full_140423305664888(0) <= fifo_full_140423305664944(1);
        
        fifo_inputs_140423305664832(0) <= outputs_140423305664888(1);
        outputs_full_140423305664888(1) <= fifo_full_140423305664832(0);
        
        fifo_inputs_140423305665000(1) <= outputs_140423305664944(0);
        outputs_full_140423305664944(0) <= fifo_full_140423305665000(1);
        
        fifo_inputs_140423305664888(0) <= outputs_140423305664944(1);
        outputs_full_140423305664944(1) <= fifo_full_140423305664888(0);
        
        fifo_inputs_140423305665056(1) <= outputs_140423305665000(0);
        outputs_full_140423305665000(0) <= fifo_full_140423305665056(1);
        
        fifo_inputs_140423305664944(0) <= outputs_140423305665000(1);
        outputs_full_140423305665000(1) <= fifo_full_140423305664944(0);
        
        fifo_inputs_140423305665112(1) <= outputs_140423305665056(0);
        outputs_full_140423305665056(0) <= fifo_full_140423305665112(1);
        
        fifo_inputs_140423305665000(0) <= outputs_140423305665056(1);
        outputs_full_140423305665056(1) <= fifo_full_140423305665000(0);
        
        fifo_inputs_140423305665168(1) <= outputs_140423305665112(0);
        outputs_full_140423305665112(0) <= fifo_full_140423305665168(1);
        
        fifo_inputs_140423305665056(0) <= outputs_140423305665112(1);
        outputs_full_140423305665112(1) <= fifo_full_140423305665056(0);
        
        fifo_inputs_140423305665224(1) <= outputs_140423305665168(0);
        outputs_full_140423305665168(0) <= fifo_full_140423305665224(1);
        
        fifo_inputs_140423305665112(0) <= outputs_140423305665168(1);
        outputs_full_140423305665168(1) <= fifo_full_140423305665112(0);
        
        fifo_inputs_140423305665280(1) <= outputs_140423305665224(0);
        outputs_full_140423305665224(0) <= fifo_full_140423305665280(1);
        
        fifo_inputs_140423305665168(0) <= outputs_140423305665224(1);
        outputs_full_140423305665224(1) <= fifo_full_140423305665168(0);
        
        fifo_inputs_140423305665336(1) <= outputs_140423305665280(0);
        outputs_full_140423305665280(0) <= fifo_full_140423305665336(1);
        
        fifo_inputs_140423305665224(0) <= outputs_140423305665280(1);
        outputs_full_140423305665280(1) <= fifo_full_140423305665224(0);
        
        fifo_inputs_140423305665392(1) <= outputs_140423305665336(0);
        outputs_full_140423305665336(0) <= fifo_full_140423305665392(1);
        
        fifo_inputs_140423305665280(0) <= outputs_140423305665336(1);
        outputs_full_140423305665336(1) <= fifo_full_140423305665280(0);
        
        fifo_inputs_140423305665448(1) <= outputs_140423305665392(0);
        outputs_full_140423305665392(0) <= fifo_full_140423305665448(1);
        
        fifo_inputs_140423305665336(0) <= outputs_140423305665392(1);
        outputs_full_140423305665392(1) <= fifo_full_140423305665336(0);
        
        fifo_inputs_140423305665504(1) <= outputs_140423305665448(0);
        outputs_full_140423305665448(0) <= fifo_full_140423305665504(1);
        
        fifo_inputs_140423305665392(0) <= outputs_140423305665448(1);
        outputs_full_140423305665448(1) <= fifo_full_140423305665392(0);
        
        fifo_inputs_140423305665560(1) <= outputs_140423305665504(0);
        outputs_full_140423305665504(0) <= fifo_full_140423305665560(1);
        
        fifo_inputs_140423305665448(0) <= outputs_140423305665504(1);
        outputs_full_140423305665504(1) <= fifo_full_140423305665448(0);
        
        fifo_inputs_140423305665616(1) <= outputs_140423305665560(0);
        outputs_full_140423305665560(0) <= fifo_full_140423305665616(1);
        
        fifo_inputs_140423305665504(0) <= outputs_140423305665560(1);
        outputs_full_140423305665560(1) <= fifo_full_140423305665504(0);
        
        fifo_inputs_140423305665672(1) <= outputs_140423305665616(0);
        outputs_full_140423305665616(0) <= fifo_full_140423305665672(1);
        
        fifo_inputs_140423305665560(0) <= outputs_140423305665616(1);
        outputs_full_140423305665616(1) <= fifo_full_140423305665560(0);
        
        fifo_inputs_140423305665728(1) <= outputs_140423305665672(0);
        outputs_full_140423305665672(0) <= fifo_full_140423305665728(1);
        
        fifo_inputs_140423305665616(0) <= outputs_140423305665672(1);
        outputs_full_140423305665672(1) <= fifo_full_140423305665616(0);
        
        fifo_inputs_140423305665784(1) <= outputs_140423305665728(0);
        outputs_full_140423305665728(0) <= fifo_full_140423305665784(1);
        
        fifo_inputs_140423305665672(0) <= outputs_140423305665728(1);
        outputs_full_140423305665728(1) <= fifo_full_140423305665672(0);
        
        fifo_inputs_140423305665840(1) <= outputs_140423305665784(0);
        outputs_full_140423305665784(0) <= fifo_full_140423305665840(1);
        
        fifo_inputs_140423305665728(0) <= outputs_140423305665784(1);
        outputs_full_140423305665784(1) <= fifo_full_140423305665728(0);
        
        fifo_inputs_140423305665896(1) <= outputs_140423305665840(0);
        outputs_full_140423305665840(0) <= fifo_full_140423305665896(1);
        
        fifo_inputs_140423305665784(0) <= outputs_140423305665840(1);
        outputs_full_140423305665840(1) <= fifo_full_140423305665784(0);
        
        fifo_inputs_140423305665952(1) <= outputs_140423305665896(0);
        outputs_full_140423305665896(0) <= fifo_full_140423305665952(1);
        
        fifo_inputs_140423305665840(0) <= outputs_140423305665896(1);
        outputs_full_140423305665896(1) <= fifo_full_140423305665840(0);
        
        fifo_inputs_140423305666008(1) <= outputs_140423305665952(0);
        outputs_full_140423305665952(0) <= fifo_full_140423305666008(1);
        
        fifo_inputs_140423305665896(0) <= outputs_140423305665952(1);
        outputs_full_140423305665952(1) <= fifo_full_140423305665896(0);
        
        fifo_inputs_140423305666064(1) <= outputs_140423305666008(0);
        outputs_full_140423305666008(0) <= fifo_full_140423305666064(1);
        
        fifo_inputs_140423305665952(0) <= outputs_140423305666008(1);
        outputs_full_140423305666008(1) <= fifo_full_140423305665952(0);
        
        fifo_inputs_140423305666120(1) <= outputs_140423305666064(0);
        outputs_full_140423305666064(0) <= fifo_full_140423305666120(1);
        
        fifo_inputs_140423305666008(0) <= outputs_140423305666064(1);
        outputs_full_140423305666064(1) <= fifo_full_140423305666008(0);
        
        fifo_inputs_140423305666176(1) <= outputs_140423305666120(0);
        outputs_full_140423305666120(0) <= fifo_full_140423305666176(1);
        
        fifo_inputs_140423305666064(0) <= outputs_140423305666120(1);
        outputs_full_140423305666120(1) <= fifo_full_140423305666064(0);
        
        fifo_inputs_140423305666232(1) <= outputs_140423305666176(0);
        outputs_full_140423305666176(0) <= fifo_full_140423305666232(1);
        
        fifo_inputs_140423305666120(0) <= outputs_140423305666176(1);
        outputs_full_140423305666176(1) <= fifo_full_140423305666120(0);
        
        fifo_inputs_140423305666288(1) <= outputs_140423305666232(0);
        outputs_full_140423305666232(0) <= fifo_full_140423305666288(1);
        
        fifo_inputs_140423305666176(0) <= outputs_140423305666232(1);
        outputs_full_140423305666232(1) <= fifo_full_140423305666176(0);
        
        fifo_inputs_140423305666344(1) <= outputs_140423305666288(0);
        outputs_full_140423305666288(0) <= fifo_full_140423305666344(1);
        
        fifo_inputs_140423305666232(0) <= outputs_140423305666288(1);
        outputs_full_140423305666288(1) <= fifo_full_140423305666232(0);
        
        fifo_inputs_140423305666400(1) <= outputs_140423305666344(0);
        outputs_full_140423305666344(0) <= fifo_full_140423305666400(1);
        
        fifo_inputs_140423305666288(0) <= outputs_140423305666344(1);
        outputs_full_140423305666344(1) <= fifo_full_140423305666288(0);
        
        fifo_inputs_140423305666456(1) <= outputs_140423305666400(0);
        outputs_full_140423305666400(0) <= fifo_full_140423305666456(1);
        
        fifo_inputs_140423305666344(0) <= outputs_140423305666400(1);
        outputs_full_140423305666400(1) <= fifo_full_140423305666344(0);
        
        fifo_inputs_140423305666512(1) <= outputs_140423305666456(0);
        outputs_full_140423305666456(0) <= fifo_full_140423305666512(1);
        
        fifo_inputs_140423305666400(0) <= outputs_140423305666456(1);
        outputs_full_140423305666456(1) <= fifo_full_140423305666400(0);
        
        fifo_inputs_140423305674824(1) <= outputs_140423305666512(0);
        outputs_full_140423305666512(0) <= fifo_full_140423305674824(1);
        
        fifo_inputs_140423305666456(0) <= outputs_140423305666512(1);
        outputs_full_140423305666512(1) <= fifo_full_140423305666456(0);
        
        fifo_inputs_140423305674880(1) <= outputs_140423305674824(0);
        outputs_full_140423305674824(0) <= fifo_full_140423305674880(1);
        
        fifo_inputs_140423305666512(0) <= outputs_140423305674824(1);
        outputs_full_140423305674824(1) <= fifo_full_140423305666512(0);
        
        fifo_inputs_140423305674936(1) <= outputs_140423305674880(0);
        outputs_full_140423305674880(0) <= fifo_full_140423305674936(1);
        
        fifo_inputs_140423305674824(0) <= outputs_140423305674880(1);
        outputs_full_140423305674880(1) <= fifo_full_140423305674824(0);
        
        fifo_inputs_140423305674992(1) <= outputs_140423305674936(0);
        outputs_full_140423305674936(0) <= fifo_full_140423305674992(1);
        
        fifo_inputs_140423305674880(0) <= outputs_140423305674936(1);
        outputs_full_140423305674936(1) <= fifo_full_140423305674880(0);
        
        fifo_inputs_140423305675048(1) <= outputs_140423305674992(0);
        outputs_full_140423305674992(0) <= fifo_full_140423305675048(1);
        
        fifo_inputs_140423305674936(0) <= outputs_140423305674992(1);
        outputs_full_140423305674992(1) <= fifo_full_140423305674936(0);
        
        fifo_inputs_140423305675104(1) <= outputs_140423305675048(0);
        outputs_full_140423305675048(0) <= fifo_full_140423305675104(1);
        
        fifo_inputs_140423305674992(0) <= outputs_140423305675048(1);
        outputs_full_140423305675048(1) <= fifo_full_140423305674992(0);
        
        fifo_inputs_140423305675160(1) <= outputs_140423305675104(0);
        outputs_full_140423305675104(0) <= fifo_full_140423305675160(1);
        
        fifo_inputs_140423305675048(0) <= outputs_140423305675104(1);
        outputs_full_140423305675104(1) <= fifo_full_140423305675048(0);
        
        fifo_inputs_140423305675216(1) <= outputs_140423305675160(0);
        outputs_full_140423305675160(0) <= fifo_full_140423305675216(1);
        
        fifo_inputs_140423305675104(0) <= outputs_140423305675160(1);
        outputs_full_140423305675160(1) <= fifo_full_140423305675104(0);
        
        fifo_inputs_140423305675272(1) <= outputs_140423305675216(0);
        outputs_full_140423305675216(0) <= fifo_full_140423305675272(1);
        
        fifo_inputs_140423305675160(0) <= outputs_140423305675216(1);
        outputs_full_140423305675216(1) <= fifo_full_140423305675160(0);
        
        fifo_inputs_140423305675328(1) <= outputs_140423305675272(0);
        outputs_full_140423305675272(0) <= fifo_full_140423305675328(1);
        
        fifo_inputs_140423305675216(0) <= outputs_140423305675272(1);
        outputs_full_140423305675272(1) <= fifo_full_140423305675216(0);
        
        fifo_inputs_140423305675384(1) <= outputs_140423305675328(0);
        outputs_full_140423305675328(0) <= fifo_full_140423305675384(1);
        
        fifo_inputs_140423305675272(0) <= outputs_140423305675328(1);
        outputs_full_140423305675328(1) <= fifo_full_140423305675272(0);
        
        fifo_inputs_140423305675440(1) <= outputs_140423305675384(0);
        outputs_full_140423305675384(0) <= fifo_full_140423305675440(1);
        
        fifo_inputs_140423305675328(0) <= outputs_140423305675384(1);
        outputs_full_140423305675384(1) <= fifo_full_140423305675328(0);
        
        fifo_inputs_140423305675496(1) <= outputs_140423305675440(0);
        outputs_full_140423305675440(0) <= fifo_full_140423305675496(1);
        
        fifo_inputs_140423305675384(0) <= outputs_140423305675440(1);
        outputs_full_140423305675440(1) <= fifo_full_140423305675384(0);
        
        fifo_inputs_140423305675552(1) <= outputs_140423305675496(0);
        outputs_full_140423305675496(0) <= fifo_full_140423305675552(1);
        
        fifo_inputs_140423305675440(0) <= outputs_140423305675496(1);
        outputs_full_140423305675496(1) <= fifo_full_140423305675440(0);
        
        fifo_inputs_140423305675608(1) <= outputs_140423305675552(0);
        outputs_full_140423305675552(0) <= fifo_full_140423305675608(1);
        
        fifo_inputs_140423305675496(0) <= outputs_140423305675552(1);
        outputs_full_140423305675552(1) <= fifo_full_140423305675496(0);
        
        fifo_inputs_140423305675664(1) <= outputs_140423305675608(0);
        outputs_full_140423305675608(0) <= fifo_full_140423305675664(1);
        
        fifo_inputs_140423305675552(0) <= outputs_140423305675608(1);
        outputs_full_140423305675608(1) <= fifo_full_140423305675552(0);
        
        fifo_inputs_140423305675720(1) <= outputs_140423305675664(0);
        outputs_full_140423305675664(0) <= fifo_full_140423305675720(1);
        
        fifo_inputs_140423305675608(0) <= outputs_140423305675664(1);
        outputs_full_140423305675664(1) <= fifo_full_140423305675608(0);
        
        fifo_inputs_140423305675664(0) <= outputs_140423305675720(1);
        outputs_full_140423305675720(1) <= fifo_full_140423305675664(0);
        

    
        core_inst_140423305571464: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305571464,
            fifo_full => fifo_full_140423305571464,
            outputs => outputs_140423305571464,
            outputs_full => outputs_full_140423305571464
        );
        
        core_inst_140423305571408: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305571408,
            fifo_full => fifo_full_140423305571408,
            outputs => outputs_140423305571408,
            outputs_full => outputs_full_140423305571408
        );
        
        core_inst_140423305571632: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305571632,
            fifo_full => fifo_full_140423305571632,
            outputs => outputs_140423305571632,
            outputs_full => outputs_full_140423305571632
        );
        
        core_inst_140423305571688: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305571688,
            fifo_full => fifo_full_140423305571688,
            outputs => outputs_140423305571688,
            outputs_full => outputs_full_140423305571688
        );
        
        core_inst_140423305571744: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305571744,
            fifo_full => fifo_full_140423305571744,
            outputs => outputs_140423305571744,
            outputs_full => outputs_full_140423305571744
        );
        
        core_inst_140423305571576: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305571576,
            fifo_full => fifo_full_140423305571576,
            outputs => outputs_140423305571576,
            outputs_full => outputs_full_140423305571576
        );
        
        core_inst_140423305571800: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305571800,
            fifo_full => fifo_full_140423305571800,
            outputs => outputs_140423305571800,
            outputs_full => outputs_full_140423305571800
        );
        
        core_inst_140423305571856: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305571856,
            fifo_full => fifo_full_140423305571856,
            outputs => outputs_140423305571856,
            outputs_full => outputs_full_140423305571856
        );
        
        core_inst_140423305571912: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305571912,
            fifo_full => fifo_full_140423305571912,
            outputs => outputs_140423305571912,
            outputs_full => outputs_full_140423305571912
        );
        
        core_inst_140423305571968: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305571968,
            fifo_full => fifo_full_140423305571968,
            outputs => outputs_140423305571968,
            outputs_full => outputs_full_140423305571968
        );
        
        core_inst_140423305571520: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305571520,
            fifo_full => fifo_full_140423305571520,
            outputs => outputs_140423305571520,
            outputs_full => outputs_full_140423305571520
        );
        
        core_inst_140423305572024: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305572024,
            fifo_full => fifo_full_140423305572024,
            outputs => outputs_140423305572024,
            outputs_full => outputs_full_140423305572024
        );
        
        core_inst_140423305572080: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305572080,
            fifo_full => fifo_full_140423305572080,
            outputs => outputs_140423305572080,
            outputs_full => outputs_full_140423305572080
        );
        
        core_inst_140423305572136: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305572136,
            fifo_full => fifo_full_140423305572136,
            outputs => outputs_140423305572136,
            outputs_full => outputs_full_140423305572136
        );
        
        core_inst_140423305572192: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305572192,
            fifo_full => fifo_full_140423305572192,
            outputs => outputs_140423305572192,
            outputs_full => outputs_full_140423305572192
        );
        
        core_inst_140423305572248: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305572248,
            fifo_full => fifo_full_140423305572248,
            outputs => outputs_140423305572248,
            outputs_full => outputs_full_140423305572248
        );
        
        core_inst_140423305572304: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305572304,
            fifo_full => fifo_full_140423305572304,
            outputs => outputs_140423305572304,
            outputs_full => outputs_full_140423305572304
        );
        
        core_inst_140423305621576: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305621576,
            fifo_full => fifo_full_140423305621576,
            outputs => outputs_140423305621576,
            outputs_full => outputs_full_140423305621576
        );
        
        core_inst_140423305621632: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305621632,
            fifo_full => fifo_full_140423305621632,
            outputs => outputs_140423305621632,
            outputs_full => outputs_full_140423305621632
        );
        
        core_inst_140423305621688: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305621688,
            fifo_full => fifo_full_140423305621688,
            outputs => outputs_140423305621688,
            outputs_full => outputs_full_140423305621688
        );
        
        core_inst_140423305621744: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305621744,
            fifo_full => fifo_full_140423305621744,
            outputs => outputs_140423305621744,
            outputs_full => outputs_full_140423305621744
        );
        
        core_inst_140423305621800: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305621800,
            fifo_full => fifo_full_140423305621800,
            outputs => outputs_140423305621800,
            outputs_full => outputs_full_140423305621800
        );
        
        core_inst_140423305621856: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305621856,
            fifo_full => fifo_full_140423305621856,
            outputs => outputs_140423305621856,
            outputs_full => outputs_full_140423305621856
        );
        
        core_inst_140423305621912: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305621912,
            fifo_full => fifo_full_140423305621912,
            outputs => outputs_140423305621912,
            outputs_full => outputs_full_140423305621912
        );
        
        core_inst_140423305621968: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305621968,
            fifo_full => fifo_full_140423305621968,
            outputs => outputs_140423305621968,
            outputs_full => outputs_full_140423305621968
        );
        
        core_inst_140423305622024: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305622024,
            fifo_full => fifo_full_140423305622024,
            outputs => outputs_140423305622024,
            outputs_full => outputs_full_140423305622024
        );
        
        core_inst_140423305622080: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305622080,
            fifo_full => fifo_full_140423305622080,
            outputs => outputs_140423305622080,
            outputs_full => outputs_full_140423305622080
        );
        
        core_inst_140423305622136: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305622136,
            fifo_full => fifo_full_140423305622136,
            outputs => outputs_140423305622136,
            outputs_full => outputs_full_140423305622136
        );
        
        core_inst_140423305622192: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305622192,
            fifo_full => fifo_full_140423305622192,
            outputs => outputs_140423305622192,
            outputs_full => outputs_full_140423305622192
        );
        
        core_inst_140423305622248: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305622248,
            fifo_full => fifo_full_140423305622248,
            outputs => outputs_140423305622248,
            outputs_full => outputs_full_140423305622248
        );
        
        core_inst_140423305622304: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305622304,
            fifo_full => fifo_full_140423305622304,
            outputs => outputs_140423305622304,
            outputs_full => outputs_full_140423305622304
        );
        
        core_inst_140423305622360: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305622360,
            fifo_full => fifo_full_140423305622360,
            outputs => outputs_140423305622360,
            outputs_full => outputs_full_140423305622360
        );
        
        core_inst_140423305622416: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305622416,
            fifo_full => fifo_full_140423305622416,
            outputs => outputs_140423305622416,
            outputs_full => outputs_full_140423305622416
        );
        
        core_inst_140423305622472: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305622472,
            fifo_full => fifo_full_140423305622472,
            outputs => outputs_140423305622472,
            outputs_full => outputs_full_140423305622472
        );
        
        core_inst_140423305622528: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305622528,
            fifo_full => fifo_full_140423305622528,
            outputs => outputs_140423305622528,
            outputs_full => outputs_full_140423305622528
        );
        
        core_inst_140423305622584: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305622584,
            fifo_full => fifo_full_140423305622584,
            outputs => outputs_140423305622584,
            outputs_full => outputs_full_140423305622584
        );
        
        core_inst_140423305622640: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305622640,
            fifo_full => fifo_full_140423305622640,
            outputs => outputs_140423305622640,
            outputs_full => outputs_full_140423305622640
        );
        
        core_inst_140423305622696: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305622696,
            fifo_full => fifo_full_140423305622696,
            outputs => outputs_140423305622696,
            outputs_full => outputs_full_140423305622696
        );
        
        core_inst_140423305622752: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305622752,
            fifo_full => fifo_full_140423305622752,
            outputs => outputs_140423305622752,
            outputs_full => outputs_full_140423305622752
        );
        
        core_inst_140423305622808: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305622808,
            fifo_full => fifo_full_140423305622808,
            outputs => outputs_140423305622808,
            outputs_full => outputs_full_140423305622808
        );
        
        core_inst_140423305622864: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305622864,
            fifo_full => fifo_full_140423305622864,
            outputs => outputs_140423305622864,
            outputs_full => outputs_full_140423305622864
        );
        
        core_inst_140423305622920: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305622920,
            fifo_full => fifo_full_140423305622920,
            outputs => outputs_140423305622920,
            outputs_full => outputs_full_140423305622920
        );
        
        core_inst_140423305622976: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305622976,
            fifo_full => fifo_full_140423305622976,
            outputs => outputs_140423305622976,
            outputs_full => outputs_full_140423305622976
        );
        
        core_inst_140423305623032: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305623032,
            fifo_full => fifo_full_140423305623032,
            outputs => outputs_140423305623032,
            outputs_full => outputs_full_140423305623032
        );
        
        core_inst_140423305623088: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305623088,
            fifo_full => fifo_full_140423305623088,
            outputs => outputs_140423305623088,
            outputs_full => outputs_full_140423305623088
        );
        
        core_inst_140423305623144: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305623144,
            fifo_full => fifo_full_140423305623144,
            outputs => outputs_140423305623144,
            outputs_full => outputs_full_140423305623144
        );
        
        core_inst_140423305623200: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305623200,
            fifo_full => fifo_full_140423305623200,
            outputs => outputs_140423305623200,
            outputs_full => outputs_full_140423305623200
        );
        
        core_inst_140423305623256: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305623256,
            fifo_full => fifo_full_140423305623256,
            outputs => outputs_140423305623256,
            outputs_full => outputs_full_140423305623256
        );
        
        core_inst_140423305623312: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305623312,
            fifo_full => fifo_full_140423305623312,
            outputs => outputs_140423305623312,
            outputs_full => outputs_full_140423305623312
        );
        
        core_inst_140423305623368: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305623368,
            fifo_full => fifo_full_140423305623368,
            outputs => outputs_140423305623368,
            outputs_full => outputs_full_140423305623368
        );
        
        core_inst_140423305623424: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305623424,
            fifo_full => fifo_full_140423305623424,
            outputs => outputs_140423305623424,
            outputs_full => outputs_full_140423305623424
        );
        
        core_inst_140423305623480: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305623480,
            fifo_full => fifo_full_140423305623480,
            outputs => outputs_140423305623480,
            outputs_full => outputs_full_140423305623480
        );
        
        core_inst_140423305623536: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305623536,
            fifo_full => fifo_full_140423305623536,
            outputs => outputs_140423305623536,
            outputs_full => outputs_full_140423305623536
        );
        
        core_inst_140423305623592: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305623592,
            fifo_full => fifo_full_140423305623592,
            outputs => outputs_140423305623592,
            outputs_full => outputs_full_140423305623592
        );
        
        core_inst_140423305623648: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305623648,
            fifo_full => fifo_full_140423305623648,
            outputs => outputs_140423305623648,
            outputs_full => outputs_full_140423305623648
        );
        
        core_inst_140423305623704: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305623704,
            fifo_full => fifo_full_140423305623704,
            outputs => outputs_140423305623704,
            outputs_full => outputs_full_140423305623704
        );
        
        core_inst_140423305623760: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305623760,
            fifo_full => fifo_full_140423305623760,
            outputs => outputs_140423305623760,
            outputs_full => outputs_full_140423305623760
        );
        
        core_inst_140423305623816: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305623816,
            fifo_full => fifo_full_140423305623816,
            outputs => outputs_140423305623816,
            outputs_full => outputs_full_140423305623816
        );
        
        core_inst_140423305623872: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305623872,
            fifo_full => fifo_full_140423305623872,
            outputs => outputs_140423305623872,
            outputs_full => outputs_full_140423305623872
        );
        
        core_inst_140423305623928: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305623928,
            fifo_full => fifo_full_140423305623928,
            outputs => outputs_140423305623928,
            outputs_full => outputs_full_140423305623928
        );
        
        core_inst_140423305623984: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305623984,
            fifo_full => fifo_full_140423305623984,
            outputs => outputs_140423305623984,
            outputs_full => outputs_full_140423305623984
        );
        
        core_inst_140423305624040: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305624040,
            fifo_full => fifo_full_140423305624040,
            outputs => outputs_140423305624040,
            outputs_full => outputs_full_140423305624040
        );
        
        core_inst_140423305624096: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305624096,
            fifo_full => fifo_full_140423305624096,
            outputs => outputs_140423305624096,
            outputs_full => outputs_full_140423305624096
        );
        
        core_inst_140423305624152: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305624152,
            fifo_full => fifo_full_140423305624152,
            outputs => outputs_140423305624152,
            outputs_full => outputs_full_140423305624152
        );
        
        core_inst_140423305624208: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305624208,
            fifo_full => fifo_full_140423305624208,
            outputs => outputs_140423305624208,
            outputs_full => outputs_full_140423305624208
        );
        
        core_inst_140423305624264: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305624264,
            fifo_full => fifo_full_140423305624264,
            outputs => outputs_140423305624264,
            outputs_full => outputs_full_140423305624264
        );
        
        core_inst_140423305624320: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305624320,
            fifo_full => fifo_full_140423305624320,
            outputs => outputs_140423305624320,
            outputs_full => outputs_full_140423305624320
        );
        
        core_inst_140423305624376: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305624376,
            fifo_full => fifo_full_140423305624376,
            outputs => outputs_140423305624376,
            outputs_full => outputs_full_140423305624376
        );
        
        core_inst_140423305624432: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305624432,
            fifo_full => fifo_full_140423305624432,
            outputs => outputs_140423305624432,
            outputs_full => outputs_full_140423305624432
        );
        
        core_inst_140423305624488: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305624488,
            fifo_full => fifo_full_140423305624488,
            outputs => outputs_140423305624488,
            outputs_full => outputs_full_140423305624488
        );
        
        core_inst_140423305624544: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305624544,
            fifo_full => fifo_full_140423305624544,
            outputs => outputs_140423305624544,
            outputs_full => outputs_full_140423305624544
        );
        
        core_inst_140423305624600: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305624600,
            fifo_full => fifo_full_140423305624600,
            outputs => outputs_140423305624600,
            outputs_full => outputs_full_140423305624600
        );
        
        core_inst_140423305624656: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305624656,
            fifo_full => fifo_full_140423305624656,
            outputs => outputs_140423305624656,
            outputs_full => outputs_full_140423305624656
        );
        
        core_inst_140423305624712: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305624712,
            fifo_full => fifo_full_140423305624712,
            outputs => outputs_140423305624712,
            outputs_full => outputs_full_140423305624712
        );
        
        core_inst_140423305624768: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305624768,
            fifo_full => fifo_full_140423305624768,
            outputs => outputs_140423305624768,
            outputs_full => outputs_full_140423305624768
        );
        
        core_inst_140423305624824: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305624824,
            fifo_full => fifo_full_140423305624824,
            outputs => outputs_140423305624824,
            outputs_full => outputs_full_140423305624824
        );
        
        core_inst_140423305624880: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305624880,
            fifo_full => fifo_full_140423305624880,
            outputs => outputs_140423305624880,
            outputs_full => outputs_full_140423305624880
        );
        
        core_inst_140423305624936: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305624936,
            fifo_full => fifo_full_140423305624936,
            outputs => outputs_140423305624936,
            outputs_full => outputs_full_140423305624936
        );
        
        core_inst_140423305624992: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305624992,
            fifo_full => fifo_full_140423305624992,
            outputs => outputs_140423305624992,
            outputs_full => outputs_full_140423305624992
        );
        
        core_inst_140423305625048: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305625048,
            fifo_full => fifo_full_140423305625048,
            outputs => outputs_140423305625048,
            outputs_full => outputs_full_140423305625048
        );
        
        core_inst_140423305625104: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305625104,
            fifo_full => fifo_full_140423305625104,
            outputs => outputs_140423305625104,
            outputs_full => outputs_full_140423305625104
        );
        
        core_inst_140423305625160: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305625160,
            fifo_full => fifo_full_140423305625160,
            outputs => outputs_140423305625160,
            outputs_full => outputs_full_140423305625160
        );
        
        core_inst_140423305625216: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305625216,
            fifo_full => fifo_full_140423305625216,
            outputs => outputs_140423305625216,
            outputs_full => outputs_full_140423305625216
        );
        
        core_inst_140423305625272: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305625272,
            fifo_full => fifo_full_140423305625272,
            outputs => outputs_140423305625272,
            outputs_full => outputs_full_140423305625272
        );
        
        core_inst_140423305625328: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305625328,
            fifo_full => fifo_full_140423305625328,
            outputs => outputs_140423305625328,
            outputs_full => outputs_full_140423305625328
        );
        
        core_inst_140423305625384: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305625384,
            fifo_full => fifo_full_140423305625384,
            outputs => outputs_140423305625384,
            outputs_full => outputs_full_140423305625384
        );
        
        core_inst_140423305625440: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305625440,
            fifo_full => fifo_full_140423305625440,
            outputs => outputs_140423305625440,
            outputs_full => outputs_full_140423305625440
        );
        
        core_inst_140423305625496: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305625496,
            fifo_full => fifo_full_140423305625496,
            outputs => outputs_140423305625496,
            outputs_full => outputs_full_140423305625496
        );
        
        core_inst_140423305625552: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305625552,
            fifo_full => fifo_full_140423305625552,
            outputs => outputs_140423305625552,
            outputs_full => outputs_full_140423305625552
        );
        
        core_inst_140423305642056: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305642056,
            fifo_full => fifo_full_140423305642056,
            outputs => outputs_140423305642056,
            outputs_full => outputs_full_140423305642056
        );
        
        core_inst_140423305642112: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305642112,
            fifo_full => fifo_full_140423305642112,
            outputs => outputs_140423305642112,
            outputs_full => outputs_full_140423305642112
        );
        
        core_inst_140423305642168: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305642168,
            fifo_full => fifo_full_140423305642168,
            outputs => outputs_140423305642168,
            outputs_full => outputs_full_140423305642168
        );
        
        core_inst_140423305642224: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305642224,
            fifo_full => fifo_full_140423305642224,
            outputs => outputs_140423305642224,
            outputs_full => outputs_full_140423305642224
        );
        
        core_inst_140423305642280: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305642280,
            fifo_full => fifo_full_140423305642280,
            outputs => outputs_140423305642280,
            outputs_full => outputs_full_140423305642280
        );
        
        core_inst_140423305642336: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305642336,
            fifo_full => fifo_full_140423305642336,
            outputs => outputs_140423305642336,
            outputs_full => outputs_full_140423305642336
        );
        
        core_inst_140423305642392: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305642392,
            fifo_full => fifo_full_140423305642392,
            outputs => outputs_140423305642392,
            outputs_full => outputs_full_140423305642392
        );
        
        core_inst_140423305642448: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305642448,
            fifo_full => fifo_full_140423305642448,
            outputs => outputs_140423305642448,
            outputs_full => outputs_full_140423305642448
        );
        
        core_inst_140423305642504: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305642504,
            fifo_full => fifo_full_140423305642504,
            outputs => outputs_140423305642504,
            outputs_full => outputs_full_140423305642504
        );
        
        core_inst_140423305642560: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305642560,
            fifo_full => fifo_full_140423305642560,
            outputs => outputs_140423305642560,
            outputs_full => outputs_full_140423305642560
        );
        
        core_inst_140423305642616: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305642616,
            fifo_full => fifo_full_140423305642616,
            outputs => outputs_140423305642616,
            outputs_full => outputs_full_140423305642616
        );
        
        core_inst_140423305642672: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305642672,
            fifo_full => fifo_full_140423305642672,
            outputs => outputs_140423305642672,
            outputs_full => outputs_full_140423305642672
        );
        
        core_inst_140423305642728: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305642728,
            fifo_full => fifo_full_140423305642728,
            outputs => outputs_140423305642728,
            outputs_full => outputs_full_140423305642728
        );
        
        core_inst_140423305642784: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305642784,
            fifo_full => fifo_full_140423305642784,
            outputs => outputs_140423305642784,
            outputs_full => outputs_full_140423305642784
        );
        
        core_inst_140423305642840: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305642840,
            fifo_full => fifo_full_140423305642840,
            outputs => outputs_140423305642840,
            outputs_full => outputs_full_140423305642840
        );
        
        core_inst_140423305642896: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305642896,
            fifo_full => fifo_full_140423305642896,
            outputs => outputs_140423305642896,
            outputs_full => outputs_full_140423305642896
        );
        
        core_inst_140423305642952: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305642952,
            fifo_full => fifo_full_140423305642952,
            outputs => outputs_140423305642952,
            outputs_full => outputs_full_140423305642952
        );
        
        core_inst_140423305643008: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305643008,
            fifo_full => fifo_full_140423305643008,
            outputs => outputs_140423305643008,
            outputs_full => outputs_full_140423305643008
        );
        
        core_inst_140423305643064: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305643064,
            fifo_full => fifo_full_140423305643064,
            outputs => outputs_140423305643064,
            outputs_full => outputs_full_140423305643064
        );
        
        core_inst_140423305643120: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305643120,
            fifo_full => fifo_full_140423305643120,
            outputs => outputs_140423305643120,
            outputs_full => outputs_full_140423305643120
        );
        
        core_inst_140423305643176: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305643176,
            fifo_full => fifo_full_140423305643176,
            outputs => outputs_140423305643176,
            outputs_full => outputs_full_140423305643176
        );
        
        core_inst_140423305643232: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305643232,
            fifo_full => fifo_full_140423305643232,
            outputs => outputs_140423305643232,
            outputs_full => outputs_full_140423305643232
        );
        
        core_inst_140423305643288: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305643288,
            fifo_full => fifo_full_140423305643288,
            outputs => outputs_140423305643288,
            outputs_full => outputs_full_140423305643288
        );
        
        core_inst_140423305643344: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305643344,
            fifo_full => fifo_full_140423305643344,
            outputs => outputs_140423305643344,
            outputs_full => outputs_full_140423305643344
        );
        
        core_inst_140423305643400: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305643400,
            fifo_full => fifo_full_140423305643400,
            outputs => outputs_140423305643400,
            outputs_full => outputs_full_140423305643400
        );
        
        core_inst_140423305643456: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305643456,
            fifo_full => fifo_full_140423305643456,
            outputs => outputs_140423305643456,
            outputs_full => outputs_full_140423305643456
        );
        
        core_inst_140423305643512: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305643512,
            fifo_full => fifo_full_140423305643512,
            outputs => outputs_140423305643512,
            outputs_full => outputs_full_140423305643512
        );
        
        core_inst_140423305643568: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305643568,
            fifo_full => fifo_full_140423305643568,
            outputs => outputs_140423305643568,
            outputs_full => outputs_full_140423305643568
        );
        
        core_inst_140423305643624: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305643624,
            fifo_full => fifo_full_140423305643624,
            outputs => outputs_140423305643624,
            outputs_full => outputs_full_140423305643624
        );
        
        core_inst_140423305643680: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305643680,
            fifo_full => fifo_full_140423305643680,
            outputs => outputs_140423305643680,
            outputs_full => outputs_full_140423305643680
        );
        
        core_inst_140423305643736: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305643736,
            fifo_full => fifo_full_140423305643736,
            outputs => outputs_140423305643736,
            outputs_full => outputs_full_140423305643736
        );
        
        core_inst_140423305643792: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305643792,
            fifo_full => fifo_full_140423305643792,
            outputs => outputs_140423305643792,
            outputs_full => outputs_full_140423305643792
        );
        
        core_inst_140423305643848: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305643848,
            fifo_full => fifo_full_140423305643848,
            outputs => outputs_140423305643848,
            outputs_full => outputs_full_140423305643848
        );
        
        core_inst_140423305643904: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305643904,
            fifo_full => fifo_full_140423305643904,
            outputs => outputs_140423305643904,
            outputs_full => outputs_full_140423305643904
        );
        
        core_inst_140423305643960: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305643960,
            fifo_full => fifo_full_140423305643960,
            outputs => outputs_140423305643960,
            outputs_full => outputs_full_140423305643960
        );
        
        core_inst_140423305644016: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305644016,
            fifo_full => fifo_full_140423305644016,
            outputs => outputs_140423305644016,
            outputs_full => outputs_full_140423305644016
        );
        
        core_inst_140423305644072: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305644072,
            fifo_full => fifo_full_140423305644072,
            outputs => outputs_140423305644072,
            outputs_full => outputs_full_140423305644072
        );
        
        core_inst_140423305644128: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305644128,
            fifo_full => fifo_full_140423305644128,
            outputs => outputs_140423305644128,
            outputs_full => outputs_full_140423305644128
        );
        
        core_inst_140423305644184: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305644184,
            fifo_full => fifo_full_140423305644184,
            outputs => outputs_140423305644184,
            outputs_full => outputs_full_140423305644184
        );
        
        core_inst_140423305644240: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305644240,
            fifo_full => fifo_full_140423305644240,
            outputs => outputs_140423305644240,
            outputs_full => outputs_full_140423305644240
        );
        
        core_inst_140423305644296: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305644296,
            fifo_full => fifo_full_140423305644296,
            outputs => outputs_140423305644296,
            outputs_full => outputs_full_140423305644296
        );
        
        core_inst_140423305644352: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305644352,
            fifo_full => fifo_full_140423305644352,
            outputs => outputs_140423305644352,
            outputs_full => outputs_full_140423305644352
        );
        
        core_inst_140423305644408: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305644408,
            fifo_full => fifo_full_140423305644408,
            outputs => outputs_140423305644408,
            outputs_full => outputs_full_140423305644408
        );
        
        core_inst_140423305644464: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305644464,
            fifo_full => fifo_full_140423305644464,
            outputs => outputs_140423305644464,
            outputs_full => outputs_full_140423305644464
        );
        
        core_inst_140423305644520: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305644520,
            fifo_full => fifo_full_140423305644520,
            outputs => outputs_140423305644520,
            outputs_full => outputs_full_140423305644520
        );
        
        core_inst_140423305644576: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305644576,
            fifo_full => fifo_full_140423305644576,
            outputs => outputs_140423305644576,
            outputs_full => outputs_full_140423305644576
        );
        
        core_inst_140423305644632: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305644632,
            fifo_full => fifo_full_140423305644632,
            outputs => outputs_140423305644632,
            outputs_full => outputs_full_140423305644632
        );
        
        core_inst_140423305644688: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305644688,
            fifo_full => fifo_full_140423305644688,
            outputs => outputs_140423305644688,
            outputs_full => outputs_full_140423305644688
        );
        
        core_inst_140423305644744: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305644744,
            fifo_full => fifo_full_140423305644744,
            outputs => outputs_140423305644744,
            outputs_full => outputs_full_140423305644744
        );
        
        core_inst_140423305644800: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305644800,
            fifo_full => fifo_full_140423305644800,
            outputs => outputs_140423305644800,
            outputs_full => outputs_full_140423305644800
        );
        
        core_inst_140423305644856: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305644856,
            fifo_full => fifo_full_140423305644856,
            outputs => outputs_140423305644856,
            outputs_full => outputs_full_140423305644856
        );
        
        core_inst_140423305644912: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305644912,
            fifo_full => fifo_full_140423305644912,
            outputs => outputs_140423305644912,
            outputs_full => outputs_full_140423305644912
        );
        
        core_inst_140423305644968: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305644968,
            fifo_full => fifo_full_140423305644968,
            outputs => outputs_140423305644968,
            outputs_full => outputs_full_140423305644968
        );
        
        core_inst_140423305645024: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305645024,
            fifo_full => fifo_full_140423305645024,
            outputs => outputs_140423305645024,
            outputs_full => outputs_full_140423305645024
        );
        
        core_inst_140423305645080: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305645080,
            fifo_full => fifo_full_140423305645080,
            outputs => outputs_140423305645080,
            outputs_full => outputs_full_140423305645080
        );
        
        core_inst_140423305645136: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305645136,
            fifo_full => fifo_full_140423305645136,
            outputs => outputs_140423305645136,
            outputs_full => outputs_full_140423305645136
        );
        
        core_inst_140423305645192: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305645192,
            fifo_full => fifo_full_140423305645192,
            outputs => outputs_140423305645192,
            outputs_full => outputs_full_140423305645192
        );
        
        core_inst_140423305645248: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305645248,
            fifo_full => fifo_full_140423305645248,
            outputs => outputs_140423305645248,
            outputs_full => outputs_full_140423305645248
        );
        
        core_inst_140423305645304: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305645304,
            fifo_full => fifo_full_140423305645304,
            outputs => outputs_140423305645304,
            outputs_full => outputs_full_140423305645304
        );
        
        core_inst_140423305645360: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305645360,
            fifo_full => fifo_full_140423305645360,
            outputs => outputs_140423305645360,
            outputs_full => outputs_full_140423305645360
        );
        
        core_inst_140423305645416: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305645416,
            fifo_full => fifo_full_140423305645416,
            outputs => outputs_140423305645416,
            outputs_full => outputs_full_140423305645416
        );
        
        core_inst_140423305645472: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305645472,
            fifo_full => fifo_full_140423305645472,
            outputs => outputs_140423305645472,
            outputs_full => outputs_full_140423305645472
        );
        
        core_inst_140423305645528: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305645528,
            fifo_full => fifo_full_140423305645528,
            outputs => outputs_140423305645528,
            outputs_full => outputs_full_140423305645528
        );
        
        core_inst_140423305645584: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305645584,
            fifo_full => fifo_full_140423305645584,
            outputs => outputs_140423305645584,
            outputs_full => outputs_full_140423305645584
        );
        
        core_inst_140423305645640: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305645640,
            fifo_full => fifo_full_140423305645640,
            outputs => outputs_140423305645640,
            outputs_full => outputs_full_140423305645640
        );
        
        core_inst_140423329706112: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423329706112,
            fifo_full => fifo_full_140423329706112,
            outputs => outputs_140423329706112,
            outputs_full => outputs_full_140423329706112
        );
        
        core_inst_140423305571240: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305571240,
            fifo_full => fifo_full_140423305571240,
            outputs => outputs_140423305571240,
            outputs_full => outputs_full_140423305571240
        );
        
        core_inst_140423305571016: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305571016,
            fifo_full => fifo_full_140423305571016,
            outputs => outputs_140423305571016,
            outputs_full => outputs_full_140423305571016
        );
        
        core_inst_140423305571296: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305571296,
            fifo_full => fifo_full_140423305571296,
            outputs => outputs_140423305571296,
            outputs_full => outputs_full_140423305571296
        );
        
        core_inst_140423305571072: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305571072,
            fifo_full => fifo_full_140423305571072,
            outputs => outputs_140423305571072,
            outputs_full => outputs_full_140423305571072
        );
        
        core_inst_140423305571128: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305571128,
            fifo_full => fifo_full_140423305571128,
            outputs => outputs_140423305571128,
            outputs_full => outputs_full_140423305571128
        );
        
        core_inst_140423305645696: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305645696,
            fifo_full => fifo_full_140423305645696,
            outputs => outputs_140423305645696,
            outputs_full => outputs_full_140423305645696
        );
        
        core_inst_140423305645752: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305645752,
            fifo_full => fifo_full_140423305645752,
            outputs => outputs_140423305645752,
            outputs_full => outputs_full_140423305645752
        );
        
        core_inst_140423305645808: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305645808,
            fifo_full => fifo_full_140423305645808,
            outputs => outputs_140423305645808,
            outputs_full => outputs_full_140423305645808
        );
        
        core_inst_140423305645864: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305645864,
            fifo_full => fifo_full_140423305645864,
            outputs => outputs_140423305645864,
            outputs_full => outputs_full_140423305645864
        );
        
        core_inst_140423305645920: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305645920,
            fifo_full => fifo_full_140423305645920,
            outputs => outputs_140423305645920,
            outputs_full => outputs_full_140423305645920
        );
        
        core_inst_140423305645976: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305645976,
            fifo_full => fifo_full_140423305645976,
            outputs => outputs_140423305645976,
            outputs_full => outputs_full_140423305645976
        );
        
        core_inst_140423305646032: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305646032,
            fifo_full => fifo_full_140423305646032,
            outputs => outputs_140423305646032,
            outputs_full => outputs_full_140423305646032
        );
        
        core_inst_140423305662536: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305662536,
            fifo_full => fifo_full_140423305662536,
            outputs => outputs_140423305662536,
            outputs_full => outputs_full_140423305662536
        );
        
        core_inst_140423305662592: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305662592,
            fifo_full => fifo_full_140423305662592,
            outputs => outputs_140423305662592,
            outputs_full => outputs_full_140423305662592
        );
        
        core_inst_140423305662648: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305662648,
            fifo_full => fifo_full_140423305662648,
            outputs => outputs_140423305662648,
            outputs_full => outputs_full_140423305662648
        );
        
        core_inst_140423305662704: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305662704,
            fifo_full => fifo_full_140423305662704,
            outputs => outputs_140423305662704,
            outputs_full => outputs_full_140423305662704
        );
        
        core_inst_140423305662760: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305662760,
            fifo_full => fifo_full_140423305662760,
            outputs => outputs_140423305662760,
            outputs_full => outputs_full_140423305662760
        );
        
        core_inst_140423305662816: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305662816,
            fifo_full => fifo_full_140423305662816,
            outputs => outputs_140423305662816,
            outputs_full => outputs_full_140423305662816
        );
        
        core_inst_140423305662872: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305662872,
            fifo_full => fifo_full_140423305662872,
            outputs => outputs_140423305662872,
            outputs_full => outputs_full_140423305662872
        );
        
        core_inst_140423305662928: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305662928,
            fifo_full => fifo_full_140423305662928,
            outputs => outputs_140423305662928,
            outputs_full => outputs_full_140423305662928
        );
        
        core_inst_140423305662984: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305662984,
            fifo_full => fifo_full_140423305662984,
            outputs => outputs_140423305662984,
            outputs_full => outputs_full_140423305662984
        );
        
        core_inst_140423305663040: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305663040,
            fifo_full => fifo_full_140423305663040,
            outputs => outputs_140423305663040,
            outputs_full => outputs_full_140423305663040
        );
        
        core_inst_140423305663096: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305663096,
            fifo_full => fifo_full_140423305663096,
            outputs => outputs_140423305663096,
            outputs_full => outputs_full_140423305663096
        );
        
        core_inst_140423305663152: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305663152,
            fifo_full => fifo_full_140423305663152,
            outputs => outputs_140423305663152,
            outputs_full => outputs_full_140423305663152
        );
        
        core_inst_140423305663208: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305663208,
            fifo_full => fifo_full_140423305663208,
            outputs => outputs_140423305663208,
            outputs_full => outputs_full_140423305663208
        );
        
        core_inst_140423305663264: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305663264,
            fifo_full => fifo_full_140423305663264,
            outputs => outputs_140423305663264,
            outputs_full => outputs_full_140423305663264
        );
        
        core_inst_140423305663320: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305663320,
            fifo_full => fifo_full_140423305663320,
            outputs => outputs_140423305663320,
            outputs_full => outputs_full_140423305663320
        );
        
        core_inst_140423305663376: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305663376,
            fifo_full => fifo_full_140423305663376,
            outputs => outputs_140423305663376,
            outputs_full => outputs_full_140423305663376
        );
        
        core_inst_140423305663432: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305663432,
            fifo_full => fifo_full_140423305663432,
            outputs => outputs_140423305663432,
            outputs_full => outputs_full_140423305663432
        );
        
        core_inst_140423305663488: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305663488,
            fifo_full => fifo_full_140423305663488,
            outputs => outputs_140423305663488,
            outputs_full => outputs_full_140423305663488
        );
        
        core_inst_140423305663544: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305663544,
            fifo_full => fifo_full_140423305663544,
            outputs => outputs_140423305663544,
            outputs_full => outputs_full_140423305663544
        );
        
        core_inst_140423305663600: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305663600,
            fifo_full => fifo_full_140423305663600,
            outputs => outputs_140423305663600,
            outputs_full => outputs_full_140423305663600
        );
        
        core_inst_140423305663656: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305663656,
            fifo_full => fifo_full_140423305663656,
            outputs => outputs_140423305663656,
            outputs_full => outputs_full_140423305663656
        );
        
        core_inst_140423305663712: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305663712,
            fifo_full => fifo_full_140423305663712,
            outputs => outputs_140423305663712,
            outputs_full => outputs_full_140423305663712
        );
        
        core_inst_140423305663768: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305663768,
            fifo_full => fifo_full_140423305663768,
            outputs => outputs_140423305663768,
            outputs_full => outputs_full_140423305663768
        );
        
        core_inst_140423305663824: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305663824,
            fifo_full => fifo_full_140423305663824,
            outputs => outputs_140423305663824,
            outputs_full => outputs_full_140423305663824
        );
        
        core_inst_140423305663880: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305663880,
            fifo_full => fifo_full_140423305663880,
            outputs => outputs_140423305663880,
            outputs_full => outputs_full_140423305663880
        );
        
        core_inst_140423305663936: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305663936,
            fifo_full => fifo_full_140423305663936,
            outputs => outputs_140423305663936,
            outputs_full => outputs_full_140423305663936
        );
        
        core_inst_140423305663992: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305663992,
            fifo_full => fifo_full_140423305663992,
            outputs => outputs_140423305663992,
            outputs_full => outputs_full_140423305663992
        );
        
        core_inst_140423305664048: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305664048,
            fifo_full => fifo_full_140423305664048,
            outputs => outputs_140423305664048,
            outputs_full => outputs_full_140423305664048
        );
        
        core_inst_140423305664104: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305664104,
            fifo_full => fifo_full_140423305664104,
            outputs => outputs_140423305664104,
            outputs_full => outputs_full_140423305664104
        );
        
        core_inst_140423305664160: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305664160,
            fifo_full => fifo_full_140423305664160,
            outputs => outputs_140423305664160,
            outputs_full => outputs_full_140423305664160
        );
        
        core_inst_140423305664216: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305664216,
            fifo_full => fifo_full_140423305664216,
            outputs => outputs_140423305664216,
            outputs_full => outputs_full_140423305664216
        );
        
        core_inst_140423305664272: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305664272,
            fifo_full => fifo_full_140423305664272,
            outputs => outputs_140423305664272,
            outputs_full => outputs_full_140423305664272
        );
        
        core_inst_140423305664328: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305664328,
            fifo_full => fifo_full_140423305664328,
            outputs => outputs_140423305664328,
            outputs_full => outputs_full_140423305664328
        );
        
        core_inst_140423305664384: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305664384,
            fifo_full => fifo_full_140423305664384,
            outputs => outputs_140423305664384,
            outputs_full => outputs_full_140423305664384
        );
        
        core_inst_140423305664440: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305664440,
            fifo_full => fifo_full_140423305664440,
            outputs => outputs_140423305664440,
            outputs_full => outputs_full_140423305664440
        );
        
        core_inst_140423305664496: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305664496,
            fifo_full => fifo_full_140423305664496,
            outputs => outputs_140423305664496,
            outputs_full => outputs_full_140423305664496
        );
        
        core_inst_140423305664552: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305664552,
            fifo_full => fifo_full_140423305664552,
            outputs => outputs_140423305664552,
            outputs_full => outputs_full_140423305664552
        );
        
        core_inst_140423305664608: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305664608,
            fifo_full => fifo_full_140423305664608,
            outputs => outputs_140423305664608,
            outputs_full => outputs_full_140423305664608
        );
        
        core_inst_140423305664664: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305664664,
            fifo_full => fifo_full_140423305664664,
            outputs => outputs_140423305664664,
            outputs_full => outputs_full_140423305664664
        );
        
        core_inst_140423305664720: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305664720,
            fifo_full => fifo_full_140423305664720,
            outputs => outputs_140423305664720,
            outputs_full => outputs_full_140423305664720
        );
        
        core_inst_140423305664776: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305664776,
            fifo_full => fifo_full_140423305664776,
            outputs => outputs_140423305664776,
            outputs_full => outputs_full_140423305664776
        );
        
        core_inst_140423305664832: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305664832,
            fifo_full => fifo_full_140423305664832,
            outputs => outputs_140423305664832,
            outputs_full => outputs_full_140423305664832
        );
        
        core_inst_140423305664888: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305664888,
            fifo_full => fifo_full_140423305664888,
            outputs => outputs_140423305664888,
            outputs_full => outputs_full_140423305664888
        );
        
        core_inst_140423305664944: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305664944,
            fifo_full => fifo_full_140423305664944,
            outputs => outputs_140423305664944,
            outputs_full => outputs_full_140423305664944
        );
        
        core_inst_140423305665000: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305665000,
            fifo_full => fifo_full_140423305665000,
            outputs => outputs_140423305665000,
            outputs_full => outputs_full_140423305665000
        );
        
        core_inst_140423305665056: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305665056,
            fifo_full => fifo_full_140423305665056,
            outputs => outputs_140423305665056,
            outputs_full => outputs_full_140423305665056
        );
        
        core_inst_140423305665112: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305665112,
            fifo_full => fifo_full_140423305665112,
            outputs => outputs_140423305665112,
            outputs_full => outputs_full_140423305665112
        );
        
        core_inst_140423305665168: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305665168,
            fifo_full => fifo_full_140423305665168,
            outputs => outputs_140423305665168,
            outputs_full => outputs_full_140423305665168
        );
        
        core_inst_140423305665224: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305665224,
            fifo_full => fifo_full_140423305665224,
            outputs => outputs_140423305665224,
            outputs_full => outputs_full_140423305665224
        );
        
        core_inst_140423305665280: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305665280,
            fifo_full => fifo_full_140423305665280,
            outputs => outputs_140423305665280,
            outputs_full => outputs_full_140423305665280
        );
        
        core_inst_140423305665336: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305665336,
            fifo_full => fifo_full_140423305665336,
            outputs => outputs_140423305665336,
            outputs_full => outputs_full_140423305665336
        );
        
        core_inst_140423305665392: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305665392,
            fifo_full => fifo_full_140423305665392,
            outputs => outputs_140423305665392,
            outputs_full => outputs_full_140423305665392
        );
        
        core_inst_140423305665448: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305665448,
            fifo_full => fifo_full_140423305665448,
            outputs => outputs_140423305665448,
            outputs_full => outputs_full_140423305665448
        );
        
        core_inst_140423305665504: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305665504,
            fifo_full => fifo_full_140423305665504,
            outputs => outputs_140423305665504,
            outputs_full => outputs_full_140423305665504
        );
        
        core_inst_140423305665560: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305665560,
            fifo_full => fifo_full_140423305665560,
            outputs => outputs_140423305665560,
            outputs_full => outputs_full_140423305665560
        );
        
        core_inst_140423305665616: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305665616,
            fifo_full => fifo_full_140423305665616,
            outputs => outputs_140423305665616,
            outputs_full => outputs_full_140423305665616
        );
        
        core_inst_140423305665672: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305665672,
            fifo_full => fifo_full_140423305665672,
            outputs => outputs_140423305665672,
            outputs_full => outputs_full_140423305665672
        );
        
        core_inst_140423305665728: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305665728,
            fifo_full => fifo_full_140423305665728,
            outputs => outputs_140423305665728,
            outputs_full => outputs_full_140423305665728
        );
        
        core_inst_140423305665784: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305665784,
            fifo_full => fifo_full_140423305665784,
            outputs => outputs_140423305665784,
            outputs_full => outputs_full_140423305665784
        );
        
        core_inst_140423305665840: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305665840,
            fifo_full => fifo_full_140423305665840,
            outputs => outputs_140423305665840,
            outputs_full => outputs_full_140423305665840
        );
        
        core_inst_140423305665896: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305665896,
            fifo_full => fifo_full_140423305665896,
            outputs => outputs_140423305665896,
            outputs_full => outputs_full_140423305665896
        );
        
        core_inst_140423305665952: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305665952,
            fifo_full => fifo_full_140423305665952,
            outputs => outputs_140423305665952,
            outputs_full => outputs_full_140423305665952
        );
        
        core_inst_140423305666008: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305666008,
            fifo_full => fifo_full_140423305666008,
            outputs => outputs_140423305666008,
            outputs_full => outputs_full_140423305666008
        );
        
        core_inst_140423305666064: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305666064,
            fifo_full => fifo_full_140423305666064,
            outputs => outputs_140423305666064,
            outputs_full => outputs_full_140423305666064
        );
        
        core_inst_140423305666120: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305666120,
            fifo_full => fifo_full_140423305666120,
            outputs => outputs_140423305666120,
            outputs_full => outputs_full_140423305666120
        );
        
        core_inst_140423305666176: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305666176,
            fifo_full => fifo_full_140423305666176,
            outputs => outputs_140423305666176,
            outputs_full => outputs_full_140423305666176
        );
        
        core_inst_140423305666232: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305666232,
            fifo_full => fifo_full_140423305666232,
            outputs => outputs_140423305666232,
            outputs_full => outputs_full_140423305666232
        );
        
        core_inst_140423305666288: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305666288,
            fifo_full => fifo_full_140423305666288,
            outputs => outputs_140423305666288,
            outputs_full => outputs_full_140423305666288
        );
        
        core_inst_140423305666344: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305666344,
            fifo_full => fifo_full_140423305666344,
            outputs => outputs_140423305666344,
            outputs_full => outputs_full_140423305666344
        );
        
        core_inst_140423305666400: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305666400,
            fifo_full => fifo_full_140423305666400,
            outputs => outputs_140423305666400,
            outputs_full => outputs_full_140423305666400
        );
        
        core_inst_140423305666456: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305666456,
            fifo_full => fifo_full_140423305666456,
            outputs => outputs_140423305666456,
            outputs_full => outputs_full_140423305666456
        );
        
        core_inst_140423305666512: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305666512,
            fifo_full => fifo_full_140423305666512,
            outputs => outputs_140423305666512,
            outputs_full => outputs_full_140423305666512
        );
        
        core_inst_140423305674824: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305674824,
            fifo_full => fifo_full_140423305674824,
            outputs => outputs_140423305674824,
            outputs_full => outputs_full_140423305674824
        );
        
        core_inst_140423305674880: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305674880,
            fifo_full => fifo_full_140423305674880,
            outputs => outputs_140423305674880,
            outputs_full => outputs_full_140423305674880
        );
        
        core_inst_140423305674936: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305674936,
            fifo_full => fifo_full_140423305674936,
            outputs => outputs_140423305674936,
            outputs_full => outputs_full_140423305674936
        );
        
        core_inst_140423305674992: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305674992,
            fifo_full => fifo_full_140423305674992,
            outputs => outputs_140423305674992,
            outputs_full => outputs_full_140423305674992
        );
        
        core_inst_140423305675048: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305675048,
            fifo_full => fifo_full_140423305675048,
            outputs => outputs_140423305675048,
            outputs_full => outputs_full_140423305675048
        );
        
        core_inst_140423305675104: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305675104,
            fifo_full => fifo_full_140423305675104,
            outputs => outputs_140423305675104,
            outputs_full => outputs_full_140423305675104
        );
        
        core_inst_140423305675160: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305675160,
            fifo_full => fifo_full_140423305675160,
            outputs => outputs_140423305675160,
            outputs_full => outputs_full_140423305675160
        );
        
        core_inst_140423305675216: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305675216,
            fifo_full => fifo_full_140423305675216,
            outputs => outputs_140423305675216,
            outputs_full => outputs_full_140423305675216
        );
        
        core_inst_140423305675272: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305675272,
            fifo_full => fifo_full_140423305675272,
            outputs => outputs_140423305675272,
            outputs_full => outputs_full_140423305675272
        );
        
        core_inst_140423305675328: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305675328,
            fifo_full => fifo_full_140423305675328,
            outputs => outputs_140423305675328,
            outputs_full => outputs_full_140423305675328
        );
        
        core_inst_140423305675384: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305675384,
            fifo_full => fifo_full_140423305675384,
            outputs => outputs_140423305675384,
            outputs_full => outputs_full_140423305675384
        );
        
        core_inst_140423305675440: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305675440,
            fifo_full => fifo_full_140423305675440,
            outputs => outputs_140423305675440,
            outputs_full => outputs_full_140423305675440
        );
        
        core_inst_140423305675496: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305675496,
            fifo_full => fifo_full_140423305675496,
            outputs => outputs_140423305675496,
            outputs_full => outputs_full_140423305675496
        );
        
        core_inst_140423305675552: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305675552,
            fifo_full => fifo_full_140423305675552,
            outputs => outputs_140423305675552,
            outputs_full => outputs_full_140423305675552
        );
        
        core_inst_140423305675608: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305675608,
            fifo_full => fifo_full_140423305675608,
            outputs => outputs_140423305675608,
            outputs_full => outputs_full_140423305675608
        );
        
        core_inst_140423305675664: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305675664,
            fifo_full => fifo_full_140423305675664,
            outputs => outputs_140423305675664,
            outputs_full => outputs_full_140423305675664
        );
        
        core_inst_140423305675720: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140423305675720,
            fifo_full => fifo_full_140423305675720,
            outputs => outputs_140423305675720,
            outputs_full => outputs_full_140423305675720
        );
        

end behav;

