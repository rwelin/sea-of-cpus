
library ieee;
use ieee.std_logic_1164.all;
use work.core_config.all;
use work.all;

entity Cube4 is
    port (
        clk: in std_logic;
        clk_en: in std_logic;
        reset: in std_logic;
        addr: in ram_addr;
        data: in word;
        we: in std_logic;
        fifo_inputs: in core_fifo_inputs_t;
        fifo_full: out std_logic_vector(0 to NUM_CORE_FIFOS-1);
        outputs: out core_fifo_inputs_t;
        outputs_full: in std_logic_vector(0 to NUM_CORE_FIFOS-1)
    );
end Cube4;

architecture behav of Cube4 is

    
        signal fifo_inputs_139730188848376: core_fifo_inputs_t;
        signal fifo_full_139730188848376: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188848376: core_fifo_inputs_t;
        signal outputs_full_139730188848376: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188848600: core_fifo_inputs_t;
        signal fifo_full_139730188848600: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188848600: core_fifo_inputs_t;
        signal outputs_full_139730188848600: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188848656: core_fifo_inputs_t;
        signal fifo_full_139730188848656: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188848656: core_fifo_inputs_t;
        signal outputs_full_139730188848656: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188848712: core_fifo_inputs_t;
        signal fifo_full_139730188848712: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188848712: core_fifo_inputs_t;
        signal outputs_full_139730188848712: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188848544: core_fifo_inputs_t;
        signal fifo_full_139730188848544: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188848544: core_fifo_inputs_t;
        signal outputs_full_139730188848544: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188848768: core_fifo_inputs_t;
        signal fifo_full_139730188848768: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188848768: core_fifo_inputs_t;
        signal outputs_full_139730188848768: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188848824: core_fifo_inputs_t;
        signal fifo_full_139730188848824: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188848824: core_fifo_inputs_t;
        signal outputs_full_139730188848824: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188848880: core_fifo_inputs_t;
        signal fifo_full_139730188848880: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188848880: core_fifo_inputs_t;
        signal outputs_full_139730188848880: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188848936: core_fifo_inputs_t;
        signal fifo_full_139730188848936: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188848936: core_fifo_inputs_t;
        signal outputs_full_139730188848936: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188848488: core_fifo_inputs_t;
        signal fifo_full_139730188848488: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188848488: core_fifo_inputs_t;
        signal outputs_full_139730188848488: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188848992: core_fifo_inputs_t;
        signal fifo_full_139730188848992: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188848992: core_fifo_inputs_t;
        signal outputs_full_139730188848992: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188849048: core_fifo_inputs_t;
        signal fifo_full_139730188849048: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188849048: core_fifo_inputs_t;
        signal outputs_full_139730188849048: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188849104: core_fifo_inputs_t;
        signal fifo_full_139730188849104: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188849104: core_fifo_inputs_t;
        signal outputs_full_139730188849104: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188894280: core_fifo_inputs_t;
        signal fifo_full_139730188894280: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188894280: core_fifo_inputs_t;
        signal outputs_full_139730188894280: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188894336: core_fifo_inputs_t;
        signal fifo_full_139730188894336: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188894336: core_fifo_inputs_t;
        signal outputs_full_139730188894336: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188894392: core_fifo_inputs_t;
        signal fifo_full_139730188894392: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188894392: core_fifo_inputs_t;
        signal outputs_full_139730188894392: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188894448: core_fifo_inputs_t;
        signal fifo_full_139730188894448: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188894448: core_fifo_inputs_t;
        signal outputs_full_139730188894448: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188894504: core_fifo_inputs_t;
        signal fifo_full_139730188894504: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188894504: core_fifo_inputs_t;
        signal outputs_full_139730188894504: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188894560: core_fifo_inputs_t;
        signal fifo_full_139730188894560: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188894560: core_fifo_inputs_t;
        signal outputs_full_139730188894560: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188894616: core_fifo_inputs_t;
        signal fifo_full_139730188894616: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188894616: core_fifo_inputs_t;
        signal outputs_full_139730188894616: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188894672: core_fifo_inputs_t;
        signal fifo_full_139730188894672: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188894672: core_fifo_inputs_t;
        signal outputs_full_139730188894672: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188894728: core_fifo_inputs_t;
        signal fifo_full_139730188894728: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188894728: core_fifo_inputs_t;
        signal outputs_full_139730188894728: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188894784: core_fifo_inputs_t;
        signal fifo_full_139730188894784: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188894784: core_fifo_inputs_t;
        signal outputs_full_139730188894784: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188894840: core_fifo_inputs_t;
        signal fifo_full_139730188894840: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188894840: core_fifo_inputs_t;
        signal outputs_full_139730188894840: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188894896: core_fifo_inputs_t;
        signal fifo_full_139730188894896: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188894896: core_fifo_inputs_t;
        signal outputs_full_139730188894896: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188894952: core_fifo_inputs_t;
        signal fifo_full_139730188894952: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188894952: core_fifo_inputs_t;
        signal outputs_full_139730188894952: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188895008: core_fifo_inputs_t;
        signal fifo_full_139730188895008: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188895008: core_fifo_inputs_t;
        signal outputs_full_139730188895008: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188895064: core_fifo_inputs_t;
        signal fifo_full_139730188895064: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188895064: core_fifo_inputs_t;
        signal outputs_full_139730188895064: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188895120: core_fifo_inputs_t;
        signal fifo_full_139730188895120: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188895120: core_fifo_inputs_t;
        signal outputs_full_139730188895120: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188895176: core_fifo_inputs_t;
        signal fifo_full_139730188895176: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188895176: core_fifo_inputs_t;
        signal outputs_full_139730188895176: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188895232: core_fifo_inputs_t;
        signal fifo_full_139730188895232: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188895232: core_fifo_inputs_t;
        signal outputs_full_139730188895232: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188895288: core_fifo_inputs_t;
        signal fifo_full_139730188895288: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188895288: core_fifo_inputs_t;
        signal outputs_full_139730188895288: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188895344: core_fifo_inputs_t;
        signal fifo_full_139730188895344: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188895344: core_fifo_inputs_t;
        signal outputs_full_139730188895344: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188895400: core_fifo_inputs_t;
        signal fifo_full_139730188895400: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188895400: core_fifo_inputs_t;
        signal outputs_full_139730188895400: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188895456: core_fifo_inputs_t;
        signal fifo_full_139730188895456: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188895456: core_fifo_inputs_t;
        signal outputs_full_139730188895456: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188895512: core_fifo_inputs_t;
        signal fifo_full_139730188895512: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188895512: core_fifo_inputs_t;
        signal outputs_full_139730188895512: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188895568: core_fifo_inputs_t;
        signal fifo_full_139730188895568: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188895568: core_fifo_inputs_t;
        signal outputs_full_139730188895568: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188895624: core_fifo_inputs_t;
        signal fifo_full_139730188895624: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188895624: core_fifo_inputs_t;
        signal outputs_full_139730188895624: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188895680: core_fifo_inputs_t;
        signal fifo_full_139730188895680: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188895680: core_fifo_inputs_t;
        signal outputs_full_139730188895680: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188895736: core_fifo_inputs_t;
        signal fifo_full_139730188895736: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188895736: core_fifo_inputs_t;
        signal outputs_full_139730188895736: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188895792: core_fifo_inputs_t;
        signal fifo_full_139730188895792: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188895792: core_fifo_inputs_t;
        signal outputs_full_139730188895792: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188895848: core_fifo_inputs_t;
        signal fifo_full_139730188895848: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188895848: core_fifo_inputs_t;
        signal outputs_full_139730188895848: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188895904: core_fifo_inputs_t;
        signal fifo_full_139730188895904: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188895904: core_fifo_inputs_t;
        signal outputs_full_139730188895904: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188895960: core_fifo_inputs_t;
        signal fifo_full_139730188895960: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188895960: core_fifo_inputs_t;
        signal outputs_full_139730188895960: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188896016: core_fifo_inputs_t;
        signal fifo_full_139730188896016: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188896016: core_fifo_inputs_t;
        signal outputs_full_139730188896016: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188896072: core_fifo_inputs_t;
        signal fifo_full_139730188896072: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188896072: core_fifo_inputs_t;
        signal outputs_full_139730188896072: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188896128: core_fifo_inputs_t;
        signal fifo_full_139730188896128: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188896128: core_fifo_inputs_t;
        signal outputs_full_139730188896128: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188896184: core_fifo_inputs_t;
        signal fifo_full_139730188896184: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188896184: core_fifo_inputs_t;
        signal outputs_full_139730188896184: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188896240: core_fifo_inputs_t;
        signal fifo_full_139730188896240: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188896240: core_fifo_inputs_t;
        signal outputs_full_139730188896240: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188896296: core_fifo_inputs_t;
        signal fifo_full_139730188896296: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188896296: core_fifo_inputs_t;
        signal outputs_full_139730188896296: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188896352: core_fifo_inputs_t;
        signal fifo_full_139730188896352: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188896352: core_fifo_inputs_t;
        signal outputs_full_139730188896352: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188896408: core_fifo_inputs_t;
        signal fifo_full_139730188896408: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188896408: core_fifo_inputs_t;
        signal outputs_full_139730188896408: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188896464: core_fifo_inputs_t;
        signal fifo_full_139730188896464: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188896464: core_fifo_inputs_t;
        signal outputs_full_139730188896464: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188896520: core_fifo_inputs_t;
        signal fifo_full_139730188896520: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188896520: core_fifo_inputs_t;
        signal outputs_full_139730188896520: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188896576: core_fifo_inputs_t;
        signal fifo_full_139730188896576: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188896576: core_fifo_inputs_t;
        signal outputs_full_139730188896576: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188896632: core_fifo_inputs_t;
        signal fifo_full_139730188896632: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188896632: core_fifo_inputs_t;
        signal outputs_full_139730188896632: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188896688: core_fifo_inputs_t;
        signal fifo_full_139730188896688: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188896688: core_fifo_inputs_t;
        signal outputs_full_139730188896688: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188896744: core_fifo_inputs_t;
        signal fifo_full_139730188896744: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188896744: core_fifo_inputs_t;
        signal outputs_full_139730188896744: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188896800: core_fifo_inputs_t;
        signal fifo_full_139730188896800: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188896800: core_fifo_inputs_t;
        signal outputs_full_139730188896800: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188896856: core_fifo_inputs_t;
        signal fifo_full_139730188896856: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188896856: core_fifo_inputs_t;
        signal outputs_full_139730188896856: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188896912: core_fifo_inputs_t;
        signal fifo_full_139730188896912: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188896912: core_fifo_inputs_t;
        signal outputs_full_139730188896912: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188896968: core_fifo_inputs_t;
        signal fifo_full_139730188896968: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188896968: core_fifo_inputs_t;
        signal outputs_full_139730188896968: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188897024: core_fifo_inputs_t;
        signal fifo_full_139730188897024: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188897024: core_fifo_inputs_t;
        signal outputs_full_139730188897024: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139730188897080: core_fifo_inputs_t;
        signal fifo_full_139730188897080: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139730188897080: core_fifo_inputs_t;
        signal outputs_full_139730188897080: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        

begin

        outputs(0) <= outputs_139730188897080(0);
        outputs_full_139730188897080(0) <= outputs_full(0);

        fifo_inputs_139730188848376(1) <= fifo_inputs(1);
        fifo_full(1) <= fifo_full_139730188848376(1);
    
        fifo_inputs_139730188848600(1) <= outputs_139730188848376(0);
        outputs_full_139730188848376(0) <= fifo_full_139730188848600(1);
        
        fifo_inputs_139730188848544(3) <= outputs_139730188848376(2);
        outputs_full_139730188848376(2) <= fifo_full_139730188848544(3);
        
        fifo_inputs_139730188894448(5) <= outputs_139730188848376(4);
        outputs_full_139730188848376(4) <= fifo_full_139730188894448(5);
        
        fifo_inputs_139730188848656(1) <= outputs_139730188848600(0);
        outputs_full_139730188848600(0) <= fifo_full_139730188848656(1);
        
        fifo_inputs_139730188848376(0) <= outputs_139730188848600(1);
        outputs_full_139730188848600(1) <= fifo_full_139730188848376(0);
        
        fifo_inputs_139730188848768(3) <= outputs_139730188848600(2);
        outputs_full_139730188848600(2) <= fifo_full_139730188848768(3);
        
        fifo_inputs_139730188894504(5) <= outputs_139730188848600(4);
        outputs_full_139730188848600(4) <= fifo_full_139730188894504(5);
        
        fifo_inputs_139730188848712(1) <= outputs_139730188848656(0);
        outputs_full_139730188848656(0) <= fifo_full_139730188848712(1);
        
        fifo_inputs_139730188848600(0) <= outputs_139730188848656(1);
        outputs_full_139730188848656(1) <= fifo_full_139730188848600(0);
        
        fifo_inputs_139730188848824(3) <= outputs_139730188848656(2);
        outputs_full_139730188848656(2) <= fifo_full_139730188848824(3);
        
        fifo_inputs_139730188894560(5) <= outputs_139730188848656(4);
        outputs_full_139730188848656(4) <= fifo_full_139730188894560(5);
        
        fifo_inputs_139730188848656(0) <= outputs_139730188848712(1);
        outputs_full_139730188848712(1) <= fifo_full_139730188848656(0);
        
        fifo_inputs_139730188848880(3) <= outputs_139730188848712(2);
        outputs_full_139730188848712(2) <= fifo_full_139730188848880(3);
        
        fifo_inputs_139730188894616(5) <= outputs_139730188848712(4);
        outputs_full_139730188848712(4) <= fifo_full_139730188894616(5);
        
        fifo_inputs_139730188848768(1) <= outputs_139730188848544(0);
        outputs_full_139730188848544(0) <= fifo_full_139730188848768(1);
        
        fifo_inputs_139730188848936(3) <= outputs_139730188848544(2);
        outputs_full_139730188848544(2) <= fifo_full_139730188848936(3);
        
        fifo_inputs_139730188848376(2) <= outputs_139730188848544(3);
        outputs_full_139730188848544(3) <= fifo_full_139730188848376(2);
        
        fifo_inputs_139730188894672(5) <= outputs_139730188848544(4);
        outputs_full_139730188848544(4) <= fifo_full_139730188894672(5);
        
        fifo_inputs_139730188848824(1) <= outputs_139730188848768(0);
        outputs_full_139730188848768(0) <= fifo_full_139730188848824(1);
        
        fifo_inputs_139730188848544(0) <= outputs_139730188848768(1);
        outputs_full_139730188848768(1) <= fifo_full_139730188848544(0);
        
        fifo_inputs_139730188848488(3) <= outputs_139730188848768(2);
        outputs_full_139730188848768(2) <= fifo_full_139730188848488(3);
        
        fifo_inputs_139730188848600(2) <= outputs_139730188848768(3);
        outputs_full_139730188848768(3) <= fifo_full_139730188848600(2);
        
        fifo_inputs_139730188894728(5) <= outputs_139730188848768(4);
        outputs_full_139730188848768(4) <= fifo_full_139730188894728(5);
        
        fifo_inputs_139730188848880(1) <= outputs_139730188848824(0);
        outputs_full_139730188848824(0) <= fifo_full_139730188848880(1);
        
        fifo_inputs_139730188848768(0) <= outputs_139730188848824(1);
        outputs_full_139730188848824(1) <= fifo_full_139730188848768(0);
        
        fifo_inputs_139730188848992(3) <= outputs_139730188848824(2);
        outputs_full_139730188848824(2) <= fifo_full_139730188848992(3);
        
        fifo_inputs_139730188848656(2) <= outputs_139730188848824(3);
        outputs_full_139730188848824(3) <= fifo_full_139730188848656(2);
        
        fifo_inputs_139730188894784(5) <= outputs_139730188848824(4);
        outputs_full_139730188848824(4) <= fifo_full_139730188894784(5);
        
        fifo_inputs_139730188848824(0) <= outputs_139730188848880(1);
        outputs_full_139730188848880(1) <= fifo_full_139730188848824(0);
        
        fifo_inputs_139730188849048(3) <= outputs_139730188848880(2);
        outputs_full_139730188848880(2) <= fifo_full_139730188849048(3);
        
        fifo_inputs_139730188848712(2) <= outputs_139730188848880(3);
        outputs_full_139730188848880(3) <= fifo_full_139730188848712(2);
        
        fifo_inputs_139730188894840(5) <= outputs_139730188848880(4);
        outputs_full_139730188848880(4) <= fifo_full_139730188894840(5);
        
        fifo_inputs_139730188848488(1) <= outputs_139730188848936(0);
        outputs_full_139730188848936(0) <= fifo_full_139730188848488(1);
        
        fifo_inputs_139730188849104(3) <= outputs_139730188848936(2);
        outputs_full_139730188848936(2) <= fifo_full_139730188849104(3);
        
        fifo_inputs_139730188848544(2) <= outputs_139730188848936(3);
        outputs_full_139730188848936(3) <= fifo_full_139730188848544(2);
        
        fifo_inputs_139730188894896(5) <= outputs_139730188848936(4);
        outputs_full_139730188848936(4) <= fifo_full_139730188894896(5);
        
        fifo_inputs_139730188848992(1) <= outputs_139730188848488(0);
        outputs_full_139730188848488(0) <= fifo_full_139730188848992(1);
        
        fifo_inputs_139730188848936(0) <= outputs_139730188848488(1);
        outputs_full_139730188848488(1) <= fifo_full_139730188848936(0);
        
        fifo_inputs_139730188894280(3) <= outputs_139730188848488(2);
        outputs_full_139730188848488(2) <= fifo_full_139730188894280(3);
        
        fifo_inputs_139730188848768(2) <= outputs_139730188848488(3);
        outputs_full_139730188848488(3) <= fifo_full_139730188848768(2);
        
        fifo_inputs_139730188894952(5) <= outputs_139730188848488(4);
        outputs_full_139730188848488(4) <= fifo_full_139730188894952(5);
        
        fifo_inputs_139730188849048(1) <= outputs_139730188848992(0);
        outputs_full_139730188848992(0) <= fifo_full_139730188849048(1);
        
        fifo_inputs_139730188848488(0) <= outputs_139730188848992(1);
        outputs_full_139730188848992(1) <= fifo_full_139730188848488(0);
        
        fifo_inputs_139730188894336(3) <= outputs_139730188848992(2);
        outputs_full_139730188848992(2) <= fifo_full_139730188894336(3);
        
        fifo_inputs_139730188848824(2) <= outputs_139730188848992(3);
        outputs_full_139730188848992(3) <= fifo_full_139730188848824(2);
        
        fifo_inputs_139730188895008(5) <= outputs_139730188848992(4);
        outputs_full_139730188848992(4) <= fifo_full_139730188895008(5);
        
        fifo_inputs_139730188848992(0) <= outputs_139730188849048(1);
        outputs_full_139730188849048(1) <= fifo_full_139730188848992(0);
        
        fifo_inputs_139730188894392(3) <= outputs_139730188849048(2);
        outputs_full_139730188849048(2) <= fifo_full_139730188894392(3);
        
        fifo_inputs_139730188848880(2) <= outputs_139730188849048(3);
        outputs_full_139730188849048(3) <= fifo_full_139730188848880(2);
        
        fifo_inputs_139730188895064(5) <= outputs_139730188849048(4);
        outputs_full_139730188849048(4) <= fifo_full_139730188895064(5);
        
        fifo_inputs_139730188894280(1) <= outputs_139730188849104(0);
        outputs_full_139730188849104(0) <= fifo_full_139730188894280(1);
        
        fifo_inputs_139730188848936(2) <= outputs_139730188849104(3);
        outputs_full_139730188849104(3) <= fifo_full_139730188848936(2);
        
        fifo_inputs_139730188895120(5) <= outputs_139730188849104(4);
        outputs_full_139730188849104(4) <= fifo_full_139730188895120(5);
        
        fifo_inputs_139730188894336(1) <= outputs_139730188894280(0);
        outputs_full_139730188894280(0) <= fifo_full_139730188894336(1);
        
        fifo_inputs_139730188849104(0) <= outputs_139730188894280(1);
        outputs_full_139730188894280(1) <= fifo_full_139730188849104(0);
        
        fifo_inputs_139730188848488(2) <= outputs_139730188894280(3);
        outputs_full_139730188894280(3) <= fifo_full_139730188848488(2);
        
        fifo_inputs_139730188895176(5) <= outputs_139730188894280(4);
        outputs_full_139730188894280(4) <= fifo_full_139730188895176(5);
        
        fifo_inputs_139730188894392(1) <= outputs_139730188894336(0);
        outputs_full_139730188894336(0) <= fifo_full_139730188894392(1);
        
        fifo_inputs_139730188894280(0) <= outputs_139730188894336(1);
        outputs_full_139730188894336(1) <= fifo_full_139730188894280(0);
        
        fifo_inputs_139730188848992(2) <= outputs_139730188894336(3);
        outputs_full_139730188894336(3) <= fifo_full_139730188848992(2);
        
        fifo_inputs_139730188895232(5) <= outputs_139730188894336(4);
        outputs_full_139730188894336(4) <= fifo_full_139730188895232(5);
        
        fifo_inputs_139730188894336(0) <= outputs_139730188894392(1);
        outputs_full_139730188894392(1) <= fifo_full_139730188894336(0);
        
        fifo_inputs_139730188849048(2) <= outputs_139730188894392(3);
        outputs_full_139730188894392(3) <= fifo_full_139730188849048(2);
        
        fifo_inputs_139730188895288(5) <= outputs_139730188894392(4);
        outputs_full_139730188894392(4) <= fifo_full_139730188895288(5);
        
        fifo_inputs_139730188894504(1) <= outputs_139730188894448(0);
        outputs_full_139730188894448(0) <= fifo_full_139730188894504(1);
        
        fifo_inputs_139730188894672(3) <= outputs_139730188894448(2);
        outputs_full_139730188894448(2) <= fifo_full_139730188894672(3);
        
        fifo_inputs_139730188895344(5) <= outputs_139730188894448(4);
        outputs_full_139730188894448(4) <= fifo_full_139730188895344(5);
        
        fifo_inputs_139730188848376(4) <= outputs_139730188894448(5);
        outputs_full_139730188894448(5) <= fifo_full_139730188848376(4);
        
        fifo_inputs_139730188894560(1) <= outputs_139730188894504(0);
        outputs_full_139730188894504(0) <= fifo_full_139730188894560(1);
        
        fifo_inputs_139730188894448(0) <= outputs_139730188894504(1);
        outputs_full_139730188894504(1) <= fifo_full_139730188894448(0);
        
        fifo_inputs_139730188894728(3) <= outputs_139730188894504(2);
        outputs_full_139730188894504(2) <= fifo_full_139730188894728(3);
        
        fifo_inputs_139730188895400(5) <= outputs_139730188894504(4);
        outputs_full_139730188894504(4) <= fifo_full_139730188895400(5);
        
        fifo_inputs_139730188848600(4) <= outputs_139730188894504(5);
        outputs_full_139730188894504(5) <= fifo_full_139730188848600(4);
        
        fifo_inputs_139730188894616(1) <= outputs_139730188894560(0);
        outputs_full_139730188894560(0) <= fifo_full_139730188894616(1);
        
        fifo_inputs_139730188894504(0) <= outputs_139730188894560(1);
        outputs_full_139730188894560(1) <= fifo_full_139730188894504(0);
        
        fifo_inputs_139730188894784(3) <= outputs_139730188894560(2);
        outputs_full_139730188894560(2) <= fifo_full_139730188894784(3);
        
        fifo_inputs_139730188895456(5) <= outputs_139730188894560(4);
        outputs_full_139730188894560(4) <= fifo_full_139730188895456(5);
        
        fifo_inputs_139730188848656(4) <= outputs_139730188894560(5);
        outputs_full_139730188894560(5) <= fifo_full_139730188848656(4);
        
        fifo_inputs_139730188894560(0) <= outputs_139730188894616(1);
        outputs_full_139730188894616(1) <= fifo_full_139730188894560(0);
        
        fifo_inputs_139730188894840(3) <= outputs_139730188894616(2);
        outputs_full_139730188894616(2) <= fifo_full_139730188894840(3);
        
        fifo_inputs_139730188895512(5) <= outputs_139730188894616(4);
        outputs_full_139730188894616(4) <= fifo_full_139730188895512(5);
        
        fifo_inputs_139730188848712(4) <= outputs_139730188894616(5);
        outputs_full_139730188894616(5) <= fifo_full_139730188848712(4);
        
        fifo_inputs_139730188894728(1) <= outputs_139730188894672(0);
        outputs_full_139730188894672(0) <= fifo_full_139730188894728(1);
        
        fifo_inputs_139730188894896(3) <= outputs_139730188894672(2);
        outputs_full_139730188894672(2) <= fifo_full_139730188894896(3);
        
        fifo_inputs_139730188894448(2) <= outputs_139730188894672(3);
        outputs_full_139730188894672(3) <= fifo_full_139730188894448(2);
        
        fifo_inputs_139730188895568(5) <= outputs_139730188894672(4);
        outputs_full_139730188894672(4) <= fifo_full_139730188895568(5);
        
        fifo_inputs_139730188848544(4) <= outputs_139730188894672(5);
        outputs_full_139730188894672(5) <= fifo_full_139730188848544(4);
        
        fifo_inputs_139730188894784(1) <= outputs_139730188894728(0);
        outputs_full_139730188894728(0) <= fifo_full_139730188894784(1);
        
        fifo_inputs_139730188894672(0) <= outputs_139730188894728(1);
        outputs_full_139730188894728(1) <= fifo_full_139730188894672(0);
        
        fifo_inputs_139730188894952(3) <= outputs_139730188894728(2);
        outputs_full_139730188894728(2) <= fifo_full_139730188894952(3);
        
        fifo_inputs_139730188894504(2) <= outputs_139730188894728(3);
        outputs_full_139730188894728(3) <= fifo_full_139730188894504(2);
        
        fifo_inputs_139730188895624(5) <= outputs_139730188894728(4);
        outputs_full_139730188894728(4) <= fifo_full_139730188895624(5);
        
        fifo_inputs_139730188848768(4) <= outputs_139730188894728(5);
        outputs_full_139730188894728(5) <= fifo_full_139730188848768(4);
        
        fifo_inputs_139730188894840(1) <= outputs_139730188894784(0);
        outputs_full_139730188894784(0) <= fifo_full_139730188894840(1);
        
        fifo_inputs_139730188894728(0) <= outputs_139730188894784(1);
        outputs_full_139730188894784(1) <= fifo_full_139730188894728(0);
        
        fifo_inputs_139730188895008(3) <= outputs_139730188894784(2);
        outputs_full_139730188894784(2) <= fifo_full_139730188895008(3);
        
        fifo_inputs_139730188894560(2) <= outputs_139730188894784(3);
        outputs_full_139730188894784(3) <= fifo_full_139730188894560(2);
        
        fifo_inputs_139730188895680(5) <= outputs_139730188894784(4);
        outputs_full_139730188894784(4) <= fifo_full_139730188895680(5);
        
        fifo_inputs_139730188848824(4) <= outputs_139730188894784(5);
        outputs_full_139730188894784(5) <= fifo_full_139730188848824(4);
        
        fifo_inputs_139730188894784(0) <= outputs_139730188894840(1);
        outputs_full_139730188894840(1) <= fifo_full_139730188894784(0);
        
        fifo_inputs_139730188895064(3) <= outputs_139730188894840(2);
        outputs_full_139730188894840(2) <= fifo_full_139730188895064(3);
        
        fifo_inputs_139730188894616(2) <= outputs_139730188894840(3);
        outputs_full_139730188894840(3) <= fifo_full_139730188894616(2);
        
        fifo_inputs_139730188895736(5) <= outputs_139730188894840(4);
        outputs_full_139730188894840(4) <= fifo_full_139730188895736(5);
        
        fifo_inputs_139730188848880(4) <= outputs_139730188894840(5);
        outputs_full_139730188894840(5) <= fifo_full_139730188848880(4);
        
        fifo_inputs_139730188894952(1) <= outputs_139730188894896(0);
        outputs_full_139730188894896(0) <= fifo_full_139730188894952(1);
        
        fifo_inputs_139730188895120(3) <= outputs_139730188894896(2);
        outputs_full_139730188894896(2) <= fifo_full_139730188895120(3);
        
        fifo_inputs_139730188894672(2) <= outputs_139730188894896(3);
        outputs_full_139730188894896(3) <= fifo_full_139730188894672(2);
        
        fifo_inputs_139730188895792(5) <= outputs_139730188894896(4);
        outputs_full_139730188894896(4) <= fifo_full_139730188895792(5);
        
        fifo_inputs_139730188848936(4) <= outputs_139730188894896(5);
        outputs_full_139730188894896(5) <= fifo_full_139730188848936(4);
        
        fifo_inputs_139730188895008(1) <= outputs_139730188894952(0);
        outputs_full_139730188894952(0) <= fifo_full_139730188895008(1);
        
        fifo_inputs_139730188894896(0) <= outputs_139730188894952(1);
        outputs_full_139730188894952(1) <= fifo_full_139730188894896(0);
        
        fifo_inputs_139730188895176(3) <= outputs_139730188894952(2);
        outputs_full_139730188894952(2) <= fifo_full_139730188895176(3);
        
        fifo_inputs_139730188894728(2) <= outputs_139730188894952(3);
        outputs_full_139730188894952(3) <= fifo_full_139730188894728(2);
        
        fifo_inputs_139730188895848(5) <= outputs_139730188894952(4);
        outputs_full_139730188894952(4) <= fifo_full_139730188895848(5);
        
        fifo_inputs_139730188848488(4) <= outputs_139730188894952(5);
        outputs_full_139730188894952(5) <= fifo_full_139730188848488(4);
        
        fifo_inputs_139730188895064(1) <= outputs_139730188895008(0);
        outputs_full_139730188895008(0) <= fifo_full_139730188895064(1);
        
        fifo_inputs_139730188894952(0) <= outputs_139730188895008(1);
        outputs_full_139730188895008(1) <= fifo_full_139730188894952(0);
        
        fifo_inputs_139730188895232(3) <= outputs_139730188895008(2);
        outputs_full_139730188895008(2) <= fifo_full_139730188895232(3);
        
        fifo_inputs_139730188894784(2) <= outputs_139730188895008(3);
        outputs_full_139730188895008(3) <= fifo_full_139730188894784(2);
        
        fifo_inputs_139730188895904(5) <= outputs_139730188895008(4);
        outputs_full_139730188895008(4) <= fifo_full_139730188895904(5);
        
        fifo_inputs_139730188848992(4) <= outputs_139730188895008(5);
        outputs_full_139730188895008(5) <= fifo_full_139730188848992(4);
        
        fifo_inputs_139730188895008(0) <= outputs_139730188895064(1);
        outputs_full_139730188895064(1) <= fifo_full_139730188895008(0);
        
        fifo_inputs_139730188895288(3) <= outputs_139730188895064(2);
        outputs_full_139730188895064(2) <= fifo_full_139730188895288(3);
        
        fifo_inputs_139730188894840(2) <= outputs_139730188895064(3);
        outputs_full_139730188895064(3) <= fifo_full_139730188894840(2);
        
        fifo_inputs_139730188895960(5) <= outputs_139730188895064(4);
        outputs_full_139730188895064(4) <= fifo_full_139730188895960(5);
        
        fifo_inputs_139730188849048(4) <= outputs_139730188895064(5);
        outputs_full_139730188895064(5) <= fifo_full_139730188849048(4);
        
        fifo_inputs_139730188895176(1) <= outputs_139730188895120(0);
        outputs_full_139730188895120(0) <= fifo_full_139730188895176(1);
        
        fifo_inputs_139730188894896(2) <= outputs_139730188895120(3);
        outputs_full_139730188895120(3) <= fifo_full_139730188894896(2);
        
        fifo_inputs_139730188896016(5) <= outputs_139730188895120(4);
        outputs_full_139730188895120(4) <= fifo_full_139730188896016(5);
        
        fifo_inputs_139730188849104(4) <= outputs_139730188895120(5);
        outputs_full_139730188895120(5) <= fifo_full_139730188849104(4);
        
        fifo_inputs_139730188895232(1) <= outputs_139730188895176(0);
        outputs_full_139730188895176(0) <= fifo_full_139730188895232(1);
        
        fifo_inputs_139730188895120(0) <= outputs_139730188895176(1);
        outputs_full_139730188895176(1) <= fifo_full_139730188895120(0);
        
        fifo_inputs_139730188894952(2) <= outputs_139730188895176(3);
        outputs_full_139730188895176(3) <= fifo_full_139730188894952(2);
        
        fifo_inputs_139730188896072(5) <= outputs_139730188895176(4);
        outputs_full_139730188895176(4) <= fifo_full_139730188896072(5);
        
        fifo_inputs_139730188894280(4) <= outputs_139730188895176(5);
        outputs_full_139730188895176(5) <= fifo_full_139730188894280(4);
        
        fifo_inputs_139730188895288(1) <= outputs_139730188895232(0);
        outputs_full_139730188895232(0) <= fifo_full_139730188895288(1);
        
        fifo_inputs_139730188895176(0) <= outputs_139730188895232(1);
        outputs_full_139730188895232(1) <= fifo_full_139730188895176(0);
        
        fifo_inputs_139730188895008(2) <= outputs_139730188895232(3);
        outputs_full_139730188895232(3) <= fifo_full_139730188895008(2);
        
        fifo_inputs_139730188896128(5) <= outputs_139730188895232(4);
        outputs_full_139730188895232(4) <= fifo_full_139730188896128(5);
        
        fifo_inputs_139730188894336(4) <= outputs_139730188895232(5);
        outputs_full_139730188895232(5) <= fifo_full_139730188894336(4);
        
        fifo_inputs_139730188895232(0) <= outputs_139730188895288(1);
        outputs_full_139730188895288(1) <= fifo_full_139730188895232(0);
        
        fifo_inputs_139730188895064(2) <= outputs_139730188895288(3);
        outputs_full_139730188895288(3) <= fifo_full_139730188895064(2);
        
        fifo_inputs_139730188896184(5) <= outputs_139730188895288(4);
        outputs_full_139730188895288(4) <= fifo_full_139730188896184(5);
        
        fifo_inputs_139730188894392(4) <= outputs_139730188895288(5);
        outputs_full_139730188895288(5) <= fifo_full_139730188894392(4);
        
        fifo_inputs_139730188895400(1) <= outputs_139730188895344(0);
        outputs_full_139730188895344(0) <= fifo_full_139730188895400(1);
        
        fifo_inputs_139730188895568(3) <= outputs_139730188895344(2);
        outputs_full_139730188895344(2) <= fifo_full_139730188895568(3);
        
        fifo_inputs_139730188896240(5) <= outputs_139730188895344(4);
        outputs_full_139730188895344(4) <= fifo_full_139730188896240(5);
        
        fifo_inputs_139730188894448(4) <= outputs_139730188895344(5);
        outputs_full_139730188895344(5) <= fifo_full_139730188894448(4);
        
        fifo_inputs_139730188895456(1) <= outputs_139730188895400(0);
        outputs_full_139730188895400(0) <= fifo_full_139730188895456(1);
        
        fifo_inputs_139730188895344(0) <= outputs_139730188895400(1);
        outputs_full_139730188895400(1) <= fifo_full_139730188895344(0);
        
        fifo_inputs_139730188895624(3) <= outputs_139730188895400(2);
        outputs_full_139730188895400(2) <= fifo_full_139730188895624(3);
        
        fifo_inputs_139730188896296(5) <= outputs_139730188895400(4);
        outputs_full_139730188895400(4) <= fifo_full_139730188896296(5);
        
        fifo_inputs_139730188894504(4) <= outputs_139730188895400(5);
        outputs_full_139730188895400(5) <= fifo_full_139730188894504(4);
        
        fifo_inputs_139730188895512(1) <= outputs_139730188895456(0);
        outputs_full_139730188895456(0) <= fifo_full_139730188895512(1);
        
        fifo_inputs_139730188895400(0) <= outputs_139730188895456(1);
        outputs_full_139730188895456(1) <= fifo_full_139730188895400(0);
        
        fifo_inputs_139730188895680(3) <= outputs_139730188895456(2);
        outputs_full_139730188895456(2) <= fifo_full_139730188895680(3);
        
        fifo_inputs_139730188896352(5) <= outputs_139730188895456(4);
        outputs_full_139730188895456(4) <= fifo_full_139730188896352(5);
        
        fifo_inputs_139730188894560(4) <= outputs_139730188895456(5);
        outputs_full_139730188895456(5) <= fifo_full_139730188894560(4);
        
        fifo_inputs_139730188895456(0) <= outputs_139730188895512(1);
        outputs_full_139730188895512(1) <= fifo_full_139730188895456(0);
        
        fifo_inputs_139730188895736(3) <= outputs_139730188895512(2);
        outputs_full_139730188895512(2) <= fifo_full_139730188895736(3);
        
        fifo_inputs_139730188896408(5) <= outputs_139730188895512(4);
        outputs_full_139730188895512(4) <= fifo_full_139730188896408(5);
        
        fifo_inputs_139730188894616(4) <= outputs_139730188895512(5);
        outputs_full_139730188895512(5) <= fifo_full_139730188894616(4);
        
        fifo_inputs_139730188895624(1) <= outputs_139730188895568(0);
        outputs_full_139730188895568(0) <= fifo_full_139730188895624(1);
        
        fifo_inputs_139730188895792(3) <= outputs_139730188895568(2);
        outputs_full_139730188895568(2) <= fifo_full_139730188895792(3);
        
        fifo_inputs_139730188895344(2) <= outputs_139730188895568(3);
        outputs_full_139730188895568(3) <= fifo_full_139730188895344(2);
        
        fifo_inputs_139730188896464(5) <= outputs_139730188895568(4);
        outputs_full_139730188895568(4) <= fifo_full_139730188896464(5);
        
        fifo_inputs_139730188894672(4) <= outputs_139730188895568(5);
        outputs_full_139730188895568(5) <= fifo_full_139730188894672(4);
        
        fifo_inputs_139730188895680(1) <= outputs_139730188895624(0);
        outputs_full_139730188895624(0) <= fifo_full_139730188895680(1);
        
        fifo_inputs_139730188895568(0) <= outputs_139730188895624(1);
        outputs_full_139730188895624(1) <= fifo_full_139730188895568(0);
        
        fifo_inputs_139730188895848(3) <= outputs_139730188895624(2);
        outputs_full_139730188895624(2) <= fifo_full_139730188895848(3);
        
        fifo_inputs_139730188895400(2) <= outputs_139730188895624(3);
        outputs_full_139730188895624(3) <= fifo_full_139730188895400(2);
        
        fifo_inputs_139730188896520(5) <= outputs_139730188895624(4);
        outputs_full_139730188895624(4) <= fifo_full_139730188896520(5);
        
        fifo_inputs_139730188894728(4) <= outputs_139730188895624(5);
        outputs_full_139730188895624(5) <= fifo_full_139730188894728(4);
        
        fifo_inputs_139730188895736(1) <= outputs_139730188895680(0);
        outputs_full_139730188895680(0) <= fifo_full_139730188895736(1);
        
        fifo_inputs_139730188895624(0) <= outputs_139730188895680(1);
        outputs_full_139730188895680(1) <= fifo_full_139730188895624(0);
        
        fifo_inputs_139730188895904(3) <= outputs_139730188895680(2);
        outputs_full_139730188895680(2) <= fifo_full_139730188895904(3);
        
        fifo_inputs_139730188895456(2) <= outputs_139730188895680(3);
        outputs_full_139730188895680(3) <= fifo_full_139730188895456(2);
        
        fifo_inputs_139730188896576(5) <= outputs_139730188895680(4);
        outputs_full_139730188895680(4) <= fifo_full_139730188896576(5);
        
        fifo_inputs_139730188894784(4) <= outputs_139730188895680(5);
        outputs_full_139730188895680(5) <= fifo_full_139730188894784(4);
        
        fifo_inputs_139730188895680(0) <= outputs_139730188895736(1);
        outputs_full_139730188895736(1) <= fifo_full_139730188895680(0);
        
        fifo_inputs_139730188895960(3) <= outputs_139730188895736(2);
        outputs_full_139730188895736(2) <= fifo_full_139730188895960(3);
        
        fifo_inputs_139730188895512(2) <= outputs_139730188895736(3);
        outputs_full_139730188895736(3) <= fifo_full_139730188895512(2);
        
        fifo_inputs_139730188896632(5) <= outputs_139730188895736(4);
        outputs_full_139730188895736(4) <= fifo_full_139730188896632(5);
        
        fifo_inputs_139730188894840(4) <= outputs_139730188895736(5);
        outputs_full_139730188895736(5) <= fifo_full_139730188894840(4);
        
        fifo_inputs_139730188895848(1) <= outputs_139730188895792(0);
        outputs_full_139730188895792(0) <= fifo_full_139730188895848(1);
        
        fifo_inputs_139730188896016(3) <= outputs_139730188895792(2);
        outputs_full_139730188895792(2) <= fifo_full_139730188896016(3);
        
        fifo_inputs_139730188895568(2) <= outputs_139730188895792(3);
        outputs_full_139730188895792(3) <= fifo_full_139730188895568(2);
        
        fifo_inputs_139730188896688(5) <= outputs_139730188895792(4);
        outputs_full_139730188895792(4) <= fifo_full_139730188896688(5);
        
        fifo_inputs_139730188894896(4) <= outputs_139730188895792(5);
        outputs_full_139730188895792(5) <= fifo_full_139730188894896(4);
        
        fifo_inputs_139730188895904(1) <= outputs_139730188895848(0);
        outputs_full_139730188895848(0) <= fifo_full_139730188895904(1);
        
        fifo_inputs_139730188895792(0) <= outputs_139730188895848(1);
        outputs_full_139730188895848(1) <= fifo_full_139730188895792(0);
        
        fifo_inputs_139730188896072(3) <= outputs_139730188895848(2);
        outputs_full_139730188895848(2) <= fifo_full_139730188896072(3);
        
        fifo_inputs_139730188895624(2) <= outputs_139730188895848(3);
        outputs_full_139730188895848(3) <= fifo_full_139730188895624(2);
        
        fifo_inputs_139730188896744(5) <= outputs_139730188895848(4);
        outputs_full_139730188895848(4) <= fifo_full_139730188896744(5);
        
        fifo_inputs_139730188894952(4) <= outputs_139730188895848(5);
        outputs_full_139730188895848(5) <= fifo_full_139730188894952(4);
        
        fifo_inputs_139730188895960(1) <= outputs_139730188895904(0);
        outputs_full_139730188895904(0) <= fifo_full_139730188895960(1);
        
        fifo_inputs_139730188895848(0) <= outputs_139730188895904(1);
        outputs_full_139730188895904(1) <= fifo_full_139730188895848(0);
        
        fifo_inputs_139730188896128(3) <= outputs_139730188895904(2);
        outputs_full_139730188895904(2) <= fifo_full_139730188896128(3);
        
        fifo_inputs_139730188895680(2) <= outputs_139730188895904(3);
        outputs_full_139730188895904(3) <= fifo_full_139730188895680(2);
        
        fifo_inputs_139730188896800(5) <= outputs_139730188895904(4);
        outputs_full_139730188895904(4) <= fifo_full_139730188896800(5);
        
        fifo_inputs_139730188895008(4) <= outputs_139730188895904(5);
        outputs_full_139730188895904(5) <= fifo_full_139730188895008(4);
        
        fifo_inputs_139730188895904(0) <= outputs_139730188895960(1);
        outputs_full_139730188895960(1) <= fifo_full_139730188895904(0);
        
        fifo_inputs_139730188896184(3) <= outputs_139730188895960(2);
        outputs_full_139730188895960(2) <= fifo_full_139730188896184(3);
        
        fifo_inputs_139730188895736(2) <= outputs_139730188895960(3);
        outputs_full_139730188895960(3) <= fifo_full_139730188895736(2);
        
        fifo_inputs_139730188896856(5) <= outputs_139730188895960(4);
        outputs_full_139730188895960(4) <= fifo_full_139730188896856(5);
        
        fifo_inputs_139730188895064(4) <= outputs_139730188895960(5);
        outputs_full_139730188895960(5) <= fifo_full_139730188895064(4);
        
        fifo_inputs_139730188896072(1) <= outputs_139730188896016(0);
        outputs_full_139730188896016(0) <= fifo_full_139730188896072(1);
        
        fifo_inputs_139730188895792(2) <= outputs_139730188896016(3);
        outputs_full_139730188896016(3) <= fifo_full_139730188895792(2);
        
        fifo_inputs_139730188896912(5) <= outputs_139730188896016(4);
        outputs_full_139730188896016(4) <= fifo_full_139730188896912(5);
        
        fifo_inputs_139730188895120(4) <= outputs_139730188896016(5);
        outputs_full_139730188896016(5) <= fifo_full_139730188895120(4);
        
        fifo_inputs_139730188896128(1) <= outputs_139730188896072(0);
        outputs_full_139730188896072(0) <= fifo_full_139730188896128(1);
        
        fifo_inputs_139730188896016(0) <= outputs_139730188896072(1);
        outputs_full_139730188896072(1) <= fifo_full_139730188896016(0);
        
        fifo_inputs_139730188895848(2) <= outputs_139730188896072(3);
        outputs_full_139730188896072(3) <= fifo_full_139730188895848(2);
        
        fifo_inputs_139730188896968(5) <= outputs_139730188896072(4);
        outputs_full_139730188896072(4) <= fifo_full_139730188896968(5);
        
        fifo_inputs_139730188895176(4) <= outputs_139730188896072(5);
        outputs_full_139730188896072(5) <= fifo_full_139730188895176(4);
        
        fifo_inputs_139730188896184(1) <= outputs_139730188896128(0);
        outputs_full_139730188896128(0) <= fifo_full_139730188896184(1);
        
        fifo_inputs_139730188896072(0) <= outputs_139730188896128(1);
        outputs_full_139730188896128(1) <= fifo_full_139730188896072(0);
        
        fifo_inputs_139730188895904(2) <= outputs_139730188896128(3);
        outputs_full_139730188896128(3) <= fifo_full_139730188895904(2);
        
        fifo_inputs_139730188897024(5) <= outputs_139730188896128(4);
        outputs_full_139730188896128(4) <= fifo_full_139730188897024(5);
        
        fifo_inputs_139730188895232(4) <= outputs_139730188896128(5);
        outputs_full_139730188896128(5) <= fifo_full_139730188895232(4);
        
        fifo_inputs_139730188896128(0) <= outputs_139730188896184(1);
        outputs_full_139730188896184(1) <= fifo_full_139730188896128(0);
        
        fifo_inputs_139730188895960(2) <= outputs_139730188896184(3);
        outputs_full_139730188896184(3) <= fifo_full_139730188895960(2);
        
        fifo_inputs_139730188897080(5) <= outputs_139730188896184(4);
        outputs_full_139730188896184(4) <= fifo_full_139730188897080(5);
        
        fifo_inputs_139730188895288(4) <= outputs_139730188896184(5);
        outputs_full_139730188896184(5) <= fifo_full_139730188895288(4);
        
        fifo_inputs_139730188896296(1) <= outputs_139730188896240(0);
        outputs_full_139730188896240(0) <= fifo_full_139730188896296(1);
        
        fifo_inputs_139730188896464(3) <= outputs_139730188896240(2);
        outputs_full_139730188896240(2) <= fifo_full_139730188896464(3);
        
        fifo_inputs_139730188895344(4) <= outputs_139730188896240(5);
        outputs_full_139730188896240(5) <= fifo_full_139730188895344(4);
        
        fifo_inputs_139730188896352(1) <= outputs_139730188896296(0);
        outputs_full_139730188896296(0) <= fifo_full_139730188896352(1);
        
        fifo_inputs_139730188896240(0) <= outputs_139730188896296(1);
        outputs_full_139730188896296(1) <= fifo_full_139730188896240(0);
        
        fifo_inputs_139730188896520(3) <= outputs_139730188896296(2);
        outputs_full_139730188896296(2) <= fifo_full_139730188896520(3);
        
        fifo_inputs_139730188895400(4) <= outputs_139730188896296(5);
        outputs_full_139730188896296(5) <= fifo_full_139730188895400(4);
        
        fifo_inputs_139730188896408(1) <= outputs_139730188896352(0);
        outputs_full_139730188896352(0) <= fifo_full_139730188896408(1);
        
        fifo_inputs_139730188896296(0) <= outputs_139730188896352(1);
        outputs_full_139730188896352(1) <= fifo_full_139730188896296(0);
        
        fifo_inputs_139730188896576(3) <= outputs_139730188896352(2);
        outputs_full_139730188896352(2) <= fifo_full_139730188896576(3);
        
        fifo_inputs_139730188895456(4) <= outputs_139730188896352(5);
        outputs_full_139730188896352(5) <= fifo_full_139730188895456(4);
        
        fifo_inputs_139730188896352(0) <= outputs_139730188896408(1);
        outputs_full_139730188896408(1) <= fifo_full_139730188896352(0);
        
        fifo_inputs_139730188896632(3) <= outputs_139730188896408(2);
        outputs_full_139730188896408(2) <= fifo_full_139730188896632(3);
        
        fifo_inputs_139730188895512(4) <= outputs_139730188896408(5);
        outputs_full_139730188896408(5) <= fifo_full_139730188895512(4);
        
        fifo_inputs_139730188896520(1) <= outputs_139730188896464(0);
        outputs_full_139730188896464(0) <= fifo_full_139730188896520(1);
        
        fifo_inputs_139730188896688(3) <= outputs_139730188896464(2);
        outputs_full_139730188896464(2) <= fifo_full_139730188896688(3);
        
        fifo_inputs_139730188896240(2) <= outputs_139730188896464(3);
        outputs_full_139730188896464(3) <= fifo_full_139730188896240(2);
        
        fifo_inputs_139730188895568(4) <= outputs_139730188896464(5);
        outputs_full_139730188896464(5) <= fifo_full_139730188895568(4);
        
        fifo_inputs_139730188896576(1) <= outputs_139730188896520(0);
        outputs_full_139730188896520(0) <= fifo_full_139730188896576(1);
        
        fifo_inputs_139730188896464(0) <= outputs_139730188896520(1);
        outputs_full_139730188896520(1) <= fifo_full_139730188896464(0);
        
        fifo_inputs_139730188896744(3) <= outputs_139730188896520(2);
        outputs_full_139730188896520(2) <= fifo_full_139730188896744(3);
        
        fifo_inputs_139730188896296(2) <= outputs_139730188896520(3);
        outputs_full_139730188896520(3) <= fifo_full_139730188896296(2);
        
        fifo_inputs_139730188895624(4) <= outputs_139730188896520(5);
        outputs_full_139730188896520(5) <= fifo_full_139730188895624(4);
        
        fifo_inputs_139730188896632(1) <= outputs_139730188896576(0);
        outputs_full_139730188896576(0) <= fifo_full_139730188896632(1);
        
        fifo_inputs_139730188896520(0) <= outputs_139730188896576(1);
        outputs_full_139730188896576(1) <= fifo_full_139730188896520(0);
        
        fifo_inputs_139730188896800(3) <= outputs_139730188896576(2);
        outputs_full_139730188896576(2) <= fifo_full_139730188896800(3);
        
        fifo_inputs_139730188896352(2) <= outputs_139730188896576(3);
        outputs_full_139730188896576(3) <= fifo_full_139730188896352(2);
        
        fifo_inputs_139730188895680(4) <= outputs_139730188896576(5);
        outputs_full_139730188896576(5) <= fifo_full_139730188895680(4);
        
        fifo_inputs_139730188896576(0) <= outputs_139730188896632(1);
        outputs_full_139730188896632(1) <= fifo_full_139730188896576(0);
        
        fifo_inputs_139730188896856(3) <= outputs_139730188896632(2);
        outputs_full_139730188896632(2) <= fifo_full_139730188896856(3);
        
        fifo_inputs_139730188896408(2) <= outputs_139730188896632(3);
        outputs_full_139730188896632(3) <= fifo_full_139730188896408(2);
        
        fifo_inputs_139730188895736(4) <= outputs_139730188896632(5);
        outputs_full_139730188896632(5) <= fifo_full_139730188895736(4);
        
        fifo_inputs_139730188896744(1) <= outputs_139730188896688(0);
        outputs_full_139730188896688(0) <= fifo_full_139730188896744(1);
        
        fifo_inputs_139730188896912(3) <= outputs_139730188896688(2);
        outputs_full_139730188896688(2) <= fifo_full_139730188896912(3);
        
        fifo_inputs_139730188896464(2) <= outputs_139730188896688(3);
        outputs_full_139730188896688(3) <= fifo_full_139730188896464(2);
        
        fifo_inputs_139730188895792(4) <= outputs_139730188896688(5);
        outputs_full_139730188896688(5) <= fifo_full_139730188895792(4);
        
        fifo_inputs_139730188896800(1) <= outputs_139730188896744(0);
        outputs_full_139730188896744(0) <= fifo_full_139730188896800(1);
        
        fifo_inputs_139730188896688(0) <= outputs_139730188896744(1);
        outputs_full_139730188896744(1) <= fifo_full_139730188896688(0);
        
        fifo_inputs_139730188896968(3) <= outputs_139730188896744(2);
        outputs_full_139730188896744(2) <= fifo_full_139730188896968(3);
        
        fifo_inputs_139730188896520(2) <= outputs_139730188896744(3);
        outputs_full_139730188896744(3) <= fifo_full_139730188896520(2);
        
        fifo_inputs_139730188895848(4) <= outputs_139730188896744(5);
        outputs_full_139730188896744(5) <= fifo_full_139730188895848(4);
        
        fifo_inputs_139730188896856(1) <= outputs_139730188896800(0);
        outputs_full_139730188896800(0) <= fifo_full_139730188896856(1);
        
        fifo_inputs_139730188896744(0) <= outputs_139730188896800(1);
        outputs_full_139730188896800(1) <= fifo_full_139730188896744(0);
        
        fifo_inputs_139730188897024(3) <= outputs_139730188896800(2);
        outputs_full_139730188896800(2) <= fifo_full_139730188897024(3);
        
        fifo_inputs_139730188896576(2) <= outputs_139730188896800(3);
        outputs_full_139730188896800(3) <= fifo_full_139730188896576(2);
        
        fifo_inputs_139730188895904(4) <= outputs_139730188896800(5);
        outputs_full_139730188896800(5) <= fifo_full_139730188895904(4);
        
        fifo_inputs_139730188896800(0) <= outputs_139730188896856(1);
        outputs_full_139730188896856(1) <= fifo_full_139730188896800(0);
        
        fifo_inputs_139730188897080(3) <= outputs_139730188896856(2);
        outputs_full_139730188896856(2) <= fifo_full_139730188897080(3);
        
        fifo_inputs_139730188896632(2) <= outputs_139730188896856(3);
        outputs_full_139730188896856(3) <= fifo_full_139730188896632(2);
        
        fifo_inputs_139730188895960(4) <= outputs_139730188896856(5);
        outputs_full_139730188896856(5) <= fifo_full_139730188895960(4);
        
        fifo_inputs_139730188896968(1) <= outputs_139730188896912(0);
        outputs_full_139730188896912(0) <= fifo_full_139730188896968(1);
        
        fifo_inputs_139730188896688(2) <= outputs_139730188896912(3);
        outputs_full_139730188896912(3) <= fifo_full_139730188896688(2);
        
        fifo_inputs_139730188896016(4) <= outputs_139730188896912(5);
        outputs_full_139730188896912(5) <= fifo_full_139730188896016(4);
        
        fifo_inputs_139730188897024(1) <= outputs_139730188896968(0);
        outputs_full_139730188896968(0) <= fifo_full_139730188897024(1);
        
        fifo_inputs_139730188896912(0) <= outputs_139730188896968(1);
        outputs_full_139730188896968(1) <= fifo_full_139730188896912(0);
        
        fifo_inputs_139730188896744(2) <= outputs_139730188896968(3);
        outputs_full_139730188896968(3) <= fifo_full_139730188896744(2);
        
        fifo_inputs_139730188896072(4) <= outputs_139730188896968(5);
        outputs_full_139730188896968(5) <= fifo_full_139730188896072(4);
        
        fifo_inputs_139730188897080(1) <= outputs_139730188897024(0);
        outputs_full_139730188897024(0) <= fifo_full_139730188897080(1);
        
        fifo_inputs_139730188896968(0) <= outputs_139730188897024(1);
        outputs_full_139730188897024(1) <= fifo_full_139730188896968(0);
        
        fifo_inputs_139730188896800(2) <= outputs_139730188897024(3);
        outputs_full_139730188897024(3) <= fifo_full_139730188896800(2);
        
        fifo_inputs_139730188896128(4) <= outputs_139730188897024(5);
        outputs_full_139730188897024(5) <= fifo_full_139730188896128(4);
        
        fifo_inputs_139730188897024(0) <= outputs_139730188897080(1);
        outputs_full_139730188897080(1) <= fifo_full_139730188897024(0);
        
        fifo_inputs_139730188896856(2) <= outputs_139730188897080(3);
        outputs_full_139730188897080(3) <= fifo_full_139730188896856(2);
        
        fifo_inputs_139730188896184(4) <= outputs_139730188897080(5);
        outputs_full_139730188897080(5) <= fifo_full_139730188896184(4);
        

    
        core_inst_139730188848376: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188848376,
            fifo_full => fifo_full_139730188848376,
            outputs => outputs_139730188848376,
            outputs_full => outputs_full_139730188848376
        );
        
        core_inst_139730188848600: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188848600,
            fifo_full => fifo_full_139730188848600,
            outputs => outputs_139730188848600,
            outputs_full => outputs_full_139730188848600
        );
        
        core_inst_139730188848656: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188848656,
            fifo_full => fifo_full_139730188848656,
            outputs => outputs_139730188848656,
            outputs_full => outputs_full_139730188848656
        );
        
        core_inst_139730188848712: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188848712,
            fifo_full => fifo_full_139730188848712,
            outputs => outputs_139730188848712,
            outputs_full => outputs_full_139730188848712
        );
        
        core_inst_139730188848544: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188848544,
            fifo_full => fifo_full_139730188848544,
            outputs => outputs_139730188848544,
            outputs_full => outputs_full_139730188848544
        );
        
        core_inst_139730188848768: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188848768,
            fifo_full => fifo_full_139730188848768,
            outputs => outputs_139730188848768,
            outputs_full => outputs_full_139730188848768
        );
        
        core_inst_139730188848824: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188848824,
            fifo_full => fifo_full_139730188848824,
            outputs => outputs_139730188848824,
            outputs_full => outputs_full_139730188848824
        );
        
        core_inst_139730188848880: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188848880,
            fifo_full => fifo_full_139730188848880,
            outputs => outputs_139730188848880,
            outputs_full => outputs_full_139730188848880
        );
        
        core_inst_139730188848936: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188848936,
            fifo_full => fifo_full_139730188848936,
            outputs => outputs_139730188848936,
            outputs_full => outputs_full_139730188848936
        );
        
        core_inst_139730188848488: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188848488,
            fifo_full => fifo_full_139730188848488,
            outputs => outputs_139730188848488,
            outputs_full => outputs_full_139730188848488
        );
        
        core_inst_139730188848992: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188848992,
            fifo_full => fifo_full_139730188848992,
            outputs => outputs_139730188848992,
            outputs_full => outputs_full_139730188848992
        );
        
        core_inst_139730188849048: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188849048,
            fifo_full => fifo_full_139730188849048,
            outputs => outputs_139730188849048,
            outputs_full => outputs_full_139730188849048
        );
        
        core_inst_139730188849104: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188849104,
            fifo_full => fifo_full_139730188849104,
            outputs => outputs_139730188849104,
            outputs_full => outputs_full_139730188849104
        );
        
        core_inst_139730188894280: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188894280,
            fifo_full => fifo_full_139730188894280,
            outputs => outputs_139730188894280,
            outputs_full => outputs_full_139730188894280
        );
        
        core_inst_139730188894336: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188894336,
            fifo_full => fifo_full_139730188894336,
            outputs => outputs_139730188894336,
            outputs_full => outputs_full_139730188894336
        );
        
        core_inst_139730188894392: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188894392,
            fifo_full => fifo_full_139730188894392,
            outputs => outputs_139730188894392,
            outputs_full => outputs_full_139730188894392
        );
        
        core_inst_139730188894448: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188894448,
            fifo_full => fifo_full_139730188894448,
            outputs => outputs_139730188894448,
            outputs_full => outputs_full_139730188894448
        );
        
        core_inst_139730188894504: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188894504,
            fifo_full => fifo_full_139730188894504,
            outputs => outputs_139730188894504,
            outputs_full => outputs_full_139730188894504
        );
        
        core_inst_139730188894560: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188894560,
            fifo_full => fifo_full_139730188894560,
            outputs => outputs_139730188894560,
            outputs_full => outputs_full_139730188894560
        );
        
        core_inst_139730188894616: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188894616,
            fifo_full => fifo_full_139730188894616,
            outputs => outputs_139730188894616,
            outputs_full => outputs_full_139730188894616
        );
        
        core_inst_139730188894672: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188894672,
            fifo_full => fifo_full_139730188894672,
            outputs => outputs_139730188894672,
            outputs_full => outputs_full_139730188894672
        );
        
        core_inst_139730188894728: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188894728,
            fifo_full => fifo_full_139730188894728,
            outputs => outputs_139730188894728,
            outputs_full => outputs_full_139730188894728
        );
        
        core_inst_139730188894784: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188894784,
            fifo_full => fifo_full_139730188894784,
            outputs => outputs_139730188894784,
            outputs_full => outputs_full_139730188894784
        );
        
        core_inst_139730188894840: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188894840,
            fifo_full => fifo_full_139730188894840,
            outputs => outputs_139730188894840,
            outputs_full => outputs_full_139730188894840
        );
        
        core_inst_139730188894896: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188894896,
            fifo_full => fifo_full_139730188894896,
            outputs => outputs_139730188894896,
            outputs_full => outputs_full_139730188894896
        );
        
        core_inst_139730188894952: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188894952,
            fifo_full => fifo_full_139730188894952,
            outputs => outputs_139730188894952,
            outputs_full => outputs_full_139730188894952
        );
        
        core_inst_139730188895008: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188895008,
            fifo_full => fifo_full_139730188895008,
            outputs => outputs_139730188895008,
            outputs_full => outputs_full_139730188895008
        );
        
        core_inst_139730188895064: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188895064,
            fifo_full => fifo_full_139730188895064,
            outputs => outputs_139730188895064,
            outputs_full => outputs_full_139730188895064
        );
        
        core_inst_139730188895120: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188895120,
            fifo_full => fifo_full_139730188895120,
            outputs => outputs_139730188895120,
            outputs_full => outputs_full_139730188895120
        );
        
        core_inst_139730188895176: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188895176,
            fifo_full => fifo_full_139730188895176,
            outputs => outputs_139730188895176,
            outputs_full => outputs_full_139730188895176
        );
        
        core_inst_139730188895232: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188895232,
            fifo_full => fifo_full_139730188895232,
            outputs => outputs_139730188895232,
            outputs_full => outputs_full_139730188895232
        );
        
        core_inst_139730188895288: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188895288,
            fifo_full => fifo_full_139730188895288,
            outputs => outputs_139730188895288,
            outputs_full => outputs_full_139730188895288
        );
        
        core_inst_139730188895344: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188895344,
            fifo_full => fifo_full_139730188895344,
            outputs => outputs_139730188895344,
            outputs_full => outputs_full_139730188895344
        );
        
        core_inst_139730188895400: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188895400,
            fifo_full => fifo_full_139730188895400,
            outputs => outputs_139730188895400,
            outputs_full => outputs_full_139730188895400
        );
        
        core_inst_139730188895456: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188895456,
            fifo_full => fifo_full_139730188895456,
            outputs => outputs_139730188895456,
            outputs_full => outputs_full_139730188895456
        );
        
        core_inst_139730188895512: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188895512,
            fifo_full => fifo_full_139730188895512,
            outputs => outputs_139730188895512,
            outputs_full => outputs_full_139730188895512
        );
        
        core_inst_139730188895568: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188895568,
            fifo_full => fifo_full_139730188895568,
            outputs => outputs_139730188895568,
            outputs_full => outputs_full_139730188895568
        );
        
        core_inst_139730188895624: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188895624,
            fifo_full => fifo_full_139730188895624,
            outputs => outputs_139730188895624,
            outputs_full => outputs_full_139730188895624
        );
        
        core_inst_139730188895680: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188895680,
            fifo_full => fifo_full_139730188895680,
            outputs => outputs_139730188895680,
            outputs_full => outputs_full_139730188895680
        );
        
        core_inst_139730188895736: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188895736,
            fifo_full => fifo_full_139730188895736,
            outputs => outputs_139730188895736,
            outputs_full => outputs_full_139730188895736
        );
        
        core_inst_139730188895792: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188895792,
            fifo_full => fifo_full_139730188895792,
            outputs => outputs_139730188895792,
            outputs_full => outputs_full_139730188895792
        );
        
        core_inst_139730188895848: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188895848,
            fifo_full => fifo_full_139730188895848,
            outputs => outputs_139730188895848,
            outputs_full => outputs_full_139730188895848
        );
        
        core_inst_139730188895904: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188895904,
            fifo_full => fifo_full_139730188895904,
            outputs => outputs_139730188895904,
            outputs_full => outputs_full_139730188895904
        );
        
        core_inst_139730188895960: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188895960,
            fifo_full => fifo_full_139730188895960,
            outputs => outputs_139730188895960,
            outputs_full => outputs_full_139730188895960
        );
        
        core_inst_139730188896016: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188896016,
            fifo_full => fifo_full_139730188896016,
            outputs => outputs_139730188896016,
            outputs_full => outputs_full_139730188896016
        );
        
        core_inst_139730188896072: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188896072,
            fifo_full => fifo_full_139730188896072,
            outputs => outputs_139730188896072,
            outputs_full => outputs_full_139730188896072
        );
        
        core_inst_139730188896128: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188896128,
            fifo_full => fifo_full_139730188896128,
            outputs => outputs_139730188896128,
            outputs_full => outputs_full_139730188896128
        );
        
        core_inst_139730188896184: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188896184,
            fifo_full => fifo_full_139730188896184,
            outputs => outputs_139730188896184,
            outputs_full => outputs_full_139730188896184
        );
        
        core_inst_139730188896240: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188896240,
            fifo_full => fifo_full_139730188896240,
            outputs => outputs_139730188896240,
            outputs_full => outputs_full_139730188896240
        );
        
        core_inst_139730188896296: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188896296,
            fifo_full => fifo_full_139730188896296,
            outputs => outputs_139730188896296,
            outputs_full => outputs_full_139730188896296
        );
        
        core_inst_139730188896352: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188896352,
            fifo_full => fifo_full_139730188896352,
            outputs => outputs_139730188896352,
            outputs_full => outputs_full_139730188896352
        );
        
        core_inst_139730188896408: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188896408,
            fifo_full => fifo_full_139730188896408,
            outputs => outputs_139730188896408,
            outputs_full => outputs_full_139730188896408
        );
        
        core_inst_139730188896464: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188896464,
            fifo_full => fifo_full_139730188896464,
            outputs => outputs_139730188896464,
            outputs_full => outputs_full_139730188896464
        );
        
        core_inst_139730188896520: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188896520,
            fifo_full => fifo_full_139730188896520,
            outputs => outputs_139730188896520,
            outputs_full => outputs_full_139730188896520
        );
        
        core_inst_139730188896576: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188896576,
            fifo_full => fifo_full_139730188896576,
            outputs => outputs_139730188896576,
            outputs_full => outputs_full_139730188896576
        );
        
        core_inst_139730188896632: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188896632,
            fifo_full => fifo_full_139730188896632,
            outputs => outputs_139730188896632,
            outputs_full => outputs_full_139730188896632
        );
        
        core_inst_139730188896688: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188896688,
            fifo_full => fifo_full_139730188896688,
            outputs => outputs_139730188896688,
            outputs_full => outputs_full_139730188896688
        );
        
        core_inst_139730188896744: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188896744,
            fifo_full => fifo_full_139730188896744,
            outputs => outputs_139730188896744,
            outputs_full => outputs_full_139730188896744
        );
        
        core_inst_139730188896800: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188896800,
            fifo_full => fifo_full_139730188896800,
            outputs => outputs_139730188896800,
            outputs_full => outputs_full_139730188896800
        );
        
        core_inst_139730188896856: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188896856,
            fifo_full => fifo_full_139730188896856,
            outputs => outputs_139730188896856,
            outputs_full => outputs_full_139730188896856
        );
        
        core_inst_139730188896912: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188896912,
            fifo_full => fifo_full_139730188896912,
            outputs => outputs_139730188896912,
            outputs_full => outputs_full_139730188896912
        );
        
        core_inst_139730188896968: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188896968,
            fifo_full => fifo_full_139730188896968,
            outputs => outputs_139730188896968,
            outputs_full => outputs_full_139730188896968
        );
        
        core_inst_139730188897024: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188897024,
            fifo_full => fifo_full_139730188897024,
            outputs => outputs_139730188897024,
            outputs_full => outputs_full_139730188897024
        );
        
        core_inst_139730188897080: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139730188897080,
            fifo_full => fifo_full_139730188897080,
            outputs => outputs_139730188897080,
            outputs_full => outputs_full_139730188897080
        );
        

end behav;

