library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity InstructionDecode is
    port (
        clk: std_logic     
    );
end InstructionDecode;

architecture behav of InstructionDecode is

begin


end behav;
