
library ieee;
use ieee.std_logic_1164.all;
use work.core_config.all;
use work.all;

entity Bichain128 is
    port (
        clk: in std_logic;
        clk_en: in std_logic;
        reset: in std_logic;
        addr: in ram_addr;
        data: in word;
        we: in std_logic;
        fifo_inputs: in core_fifo_inputs_t;
        fifo_full: out std_logic_vector(0 to NUM_CORE_FIFOS-1);
        outputs: out core_fifo_inputs_t;
        outputs_full: in std_logic_vector(0 to NUM_CORE_FIFOS-1)
    );
end Bichain128;

architecture behav of Bichain128 is

    
        signal fifo_inputs_140248006679688: core_fifo_inputs_t;
        signal fifo_full_140248006679688: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006679688: core_fifo_inputs_t;
        signal outputs_full_140248006679688: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006679632: core_fifo_inputs_t;
        signal fifo_full_140248006679632: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006679632: core_fifo_inputs_t;
        signal outputs_full_140248006679632: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006679856: core_fifo_inputs_t;
        signal fifo_full_140248006679856: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006679856: core_fifo_inputs_t;
        signal outputs_full_140248006679856: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006679912: core_fifo_inputs_t;
        signal fifo_full_140248006679912: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006679912: core_fifo_inputs_t;
        signal outputs_full_140248006679912: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006679968: core_fifo_inputs_t;
        signal fifo_full_140248006679968: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006679968: core_fifo_inputs_t;
        signal outputs_full_140248006679968: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006679800: core_fifo_inputs_t;
        signal fifo_full_140248006679800: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006679800: core_fifo_inputs_t;
        signal outputs_full_140248006679800: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006680024: core_fifo_inputs_t;
        signal fifo_full_140248006680024: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006680024: core_fifo_inputs_t;
        signal outputs_full_140248006680024: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006680080: core_fifo_inputs_t;
        signal fifo_full_140248006680080: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006680080: core_fifo_inputs_t;
        signal outputs_full_140248006680080: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006680136: core_fifo_inputs_t;
        signal fifo_full_140248006680136: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006680136: core_fifo_inputs_t;
        signal outputs_full_140248006680136: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006680192: core_fifo_inputs_t;
        signal fifo_full_140248006680192: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006680192: core_fifo_inputs_t;
        signal outputs_full_140248006680192: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006679744: core_fifo_inputs_t;
        signal fifo_full_140248006679744: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006679744: core_fifo_inputs_t;
        signal outputs_full_140248006679744: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006680248: core_fifo_inputs_t;
        signal fifo_full_140248006680248: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006680248: core_fifo_inputs_t;
        signal outputs_full_140248006680248: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006680304: core_fifo_inputs_t;
        signal fifo_full_140248006680304: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006680304: core_fifo_inputs_t;
        signal outputs_full_140248006680304: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006680360: core_fifo_inputs_t;
        signal fifo_full_140248006680360: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006680360: core_fifo_inputs_t;
        signal outputs_full_140248006680360: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006680416: core_fifo_inputs_t;
        signal fifo_full_140248006680416: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006680416: core_fifo_inputs_t;
        signal outputs_full_140248006680416: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006680472: core_fifo_inputs_t;
        signal fifo_full_140248006680472: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006680472: core_fifo_inputs_t;
        signal outputs_full_140248006680472: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006680528: core_fifo_inputs_t;
        signal fifo_full_140248006680528: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006680528: core_fifo_inputs_t;
        signal outputs_full_140248006680528: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006729800: core_fifo_inputs_t;
        signal fifo_full_140248006729800: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006729800: core_fifo_inputs_t;
        signal outputs_full_140248006729800: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006729856: core_fifo_inputs_t;
        signal fifo_full_140248006729856: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006729856: core_fifo_inputs_t;
        signal outputs_full_140248006729856: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006729912: core_fifo_inputs_t;
        signal fifo_full_140248006729912: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006729912: core_fifo_inputs_t;
        signal outputs_full_140248006729912: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006729968: core_fifo_inputs_t;
        signal fifo_full_140248006729968: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006729968: core_fifo_inputs_t;
        signal outputs_full_140248006729968: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006730024: core_fifo_inputs_t;
        signal fifo_full_140248006730024: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006730024: core_fifo_inputs_t;
        signal outputs_full_140248006730024: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006730080: core_fifo_inputs_t;
        signal fifo_full_140248006730080: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006730080: core_fifo_inputs_t;
        signal outputs_full_140248006730080: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006730136: core_fifo_inputs_t;
        signal fifo_full_140248006730136: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006730136: core_fifo_inputs_t;
        signal outputs_full_140248006730136: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006730192: core_fifo_inputs_t;
        signal fifo_full_140248006730192: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006730192: core_fifo_inputs_t;
        signal outputs_full_140248006730192: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006730248: core_fifo_inputs_t;
        signal fifo_full_140248006730248: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006730248: core_fifo_inputs_t;
        signal outputs_full_140248006730248: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006730304: core_fifo_inputs_t;
        signal fifo_full_140248006730304: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006730304: core_fifo_inputs_t;
        signal outputs_full_140248006730304: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006730360: core_fifo_inputs_t;
        signal fifo_full_140248006730360: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006730360: core_fifo_inputs_t;
        signal outputs_full_140248006730360: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006730416: core_fifo_inputs_t;
        signal fifo_full_140248006730416: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006730416: core_fifo_inputs_t;
        signal outputs_full_140248006730416: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006730472: core_fifo_inputs_t;
        signal fifo_full_140248006730472: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006730472: core_fifo_inputs_t;
        signal outputs_full_140248006730472: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006730528: core_fifo_inputs_t;
        signal fifo_full_140248006730528: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006730528: core_fifo_inputs_t;
        signal outputs_full_140248006730528: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006730584: core_fifo_inputs_t;
        signal fifo_full_140248006730584: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006730584: core_fifo_inputs_t;
        signal outputs_full_140248006730584: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006730640: core_fifo_inputs_t;
        signal fifo_full_140248006730640: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006730640: core_fifo_inputs_t;
        signal outputs_full_140248006730640: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006730696: core_fifo_inputs_t;
        signal fifo_full_140248006730696: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006730696: core_fifo_inputs_t;
        signal outputs_full_140248006730696: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006730752: core_fifo_inputs_t;
        signal fifo_full_140248006730752: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006730752: core_fifo_inputs_t;
        signal outputs_full_140248006730752: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006730808: core_fifo_inputs_t;
        signal fifo_full_140248006730808: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006730808: core_fifo_inputs_t;
        signal outputs_full_140248006730808: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006730864: core_fifo_inputs_t;
        signal fifo_full_140248006730864: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006730864: core_fifo_inputs_t;
        signal outputs_full_140248006730864: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006730920: core_fifo_inputs_t;
        signal fifo_full_140248006730920: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006730920: core_fifo_inputs_t;
        signal outputs_full_140248006730920: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006730976: core_fifo_inputs_t;
        signal fifo_full_140248006730976: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006730976: core_fifo_inputs_t;
        signal outputs_full_140248006730976: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006731032: core_fifo_inputs_t;
        signal fifo_full_140248006731032: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006731032: core_fifo_inputs_t;
        signal outputs_full_140248006731032: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006731088: core_fifo_inputs_t;
        signal fifo_full_140248006731088: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006731088: core_fifo_inputs_t;
        signal outputs_full_140248006731088: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006731144: core_fifo_inputs_t;
        signal fifo_full_140248006731144: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006731144: core_fifo_inputs_t;
        signal outputs_full_140248006731144: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006731200: core_fifo_inputs_t;
        signal fifo_full_140248006731200: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006731200: core_fifo_inputs_t;
        signal outputs_full_140248006731200: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006731256: core_fifo_inputs_t;
        signal fifo_full_140248006731256: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006731256: core_fifo_inputs_t;
        signal outputs_full_140248006731256: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006731312: core_fifo_inputs_t;
        signal fifo_full_140248006731312: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006731312: core_fifo_inputs_t;
        signal outputs_full_140248006731312: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006731368: core_fifo_inputs_t;
        signal fifo_full_140248006731368: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006731368: core_fifo_inputs_t;
        signal outputs_full_140248006731368: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006731424: core_fifo_inputs_t;
        signal fifo_full_140248006731424: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006731424: core_fifo_inputs_t;
        signal outputs_full_140248006731424: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006731480: core_fifo_inputs_t;
        signal fifo_full_140248006731480: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006731480: core_fifo_inputs_t;
        signal outputs_full_140248006731480: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006731536: core_fifo_inputs_t;
        signal fifo_full_140248006731536: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006731536: core_fifo_inputs_t;
        signal outputs_full_140248006731536: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006731592: core_fifo_inputs_t;
        signal fifo_full_140248006731592: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006731592: core_fifo_inputs_t;
        signal outputs_full_140248006731592: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006731648: core_fifo_inputs_t;
        signal fifo_full_140248006731648: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006731648: core_fifo_inputs_t;
        signal outputs_full_140248006731648: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006731704: core_fifo_inputs_t;
        signal fifo_full_140248006731704: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006731704: core_fifo_inputs_t;
        signal outputs_full_140248006731704: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006731760: core_fifo_inputs_t;
        signal fifo_full_140248006731760: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006731760: core_fifo_inputs_t;
        signal outputs_full_140248006731760: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006731816: core_fifo_inputs_t;
        signal fifo_full_140248006731816: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006731816: core_fifo_inputs_t;
        signal outputs_full_140248006731816: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006731872: core_fifo_inputs_t;
        signal fifo_full_140248006731872: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006731872: core_fifo_inputs_t;
        signal outputs_full_140248006731872: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006731928: core_fifo_inputs_t;
        signal fifo_full_140248006731928: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006731928: core_fifo_inputs_t;
        signal outputs_full_140248006731928: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006731984: core_fifo_inputs_t;
        signal fifo_full_140248006731984: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006731984: core_fifo_inputs_t;
        signal outputs_full_140248006731984: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006732040: core_fifo_inputs_t;
        signal fifo_full_140248006732040: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006732040: core_fifo_inputs_t;
        signal outputs_full_140248006732040: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006732096: core_fifo_inputs_t;
        signal fifo_full_140248006732096: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006732096: core_fifo_inputs_t;
        signal outputs_full_140248006732096: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006732152: core_fifo_inputs_t;
        signal fifo_full_140248006732152: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006732152: core_fifo_inputs_t;
        signal outputs_full_140248006732152: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006732208: core_fifo_inputs_t;
        signal fifo_full_140248006732208: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006732208: core_fifo_inputs_t;
        signal outputs_full_140248006732208: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006732264: core_fifo_inputs_t;
        signal fifo_full_140248006732264: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006732264: core_fifo_inputs_t;
        signal outputs_full_140248006732264: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006732320: core_fifo_inputs_t;
        signal fifo_full_140248006732320: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006732320: core_fifo_inputs_t;
        signal outputs_full_140248006732320: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006732376: core_fifo_inputs_t;
        signal fifo_full_140248006732376: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006732376: core_fifo_inputs_t;
        signal outputs_full_140248006732376: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006732432: core_fifo_inputs_t;
        signal fifo_full_140248006732432: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006732432: core_fifo_inputs_t;
        signal outputs_full_140248006732432: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006732488: core_fifo_inputs_t;
        signal fifo_full_140248006732488: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006732488: core_fifo_inputs_t;
        signal outputs_full_140248006732488: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006732544: core_fifo_inputs_t;
        signal fifo_full_140248006732544: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006732544: core_fifo_inputs_t;
        signal outputs_full_140248006732544: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006732600: core_fifo_inputs_t;
        signal fifo_full_140248006732600: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006732600: core_fifo_inputs_t;
        signal outputs_full_140248006732600: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006732656: core_fifo_inputs_t;
        signal fifo_full_140248006732656: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006732656: core_fifo_inputs_t;
        signal outputs_full_140248006732656: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006732712: core_fifo_inputs_t;
        signal fifo_full_140248006732712: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006732712: core_fifo_inputs_t;
        signal outputs_full_140248006732712: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006732768: core_fifo_inputs_t;
        signal fifo_full_140248006732768: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006732768: core_fifo_inputs_t;
        signal outputs_full_140248006732768: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006732824: core_fifo_inputs_t;
        signal fifo_full_140248006732824: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006732824: core_fifo_inputs_t;
        signal outputs_full_140248006732824: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006732880: core_fifo_inputs_t;
        signal fifo_full_140248006732880: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006732880: core_fifo_inputs_t;
        signal outputs_full_140248006732880: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006732936: core_fifo_inputs_t;
        signal fifo_full_140248006732936: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006732936: core_fifo_inputs_t;
        signal outputs_full_140248006732936: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006732992: core_fifo_inputs_t;
        signal fifo_full_140248006732992: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006732992: core_fifo_inputs_t;
        signal outputs_full_140248006732992: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006733048: core_fifo_inputs_t;
        signal fifo_full_140248006733048: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006733048: core_fifo_inputs_t;
        signal outputs_full_140248006733048: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006733104: core_fifo_inputs_t;
        signal fifo_full_140248006733104: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006733104: core_fifo_inputs_t;
        signal outputs_full_140248006733104: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006733160: core_fifo_inputs_t;
        signal fifo_full_140248006733160: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006733160: core_fifo_inputs_t;
        signal outputs_full_140248006733160: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006733216: core_fifo_inputs_t;
        signal fifo_full_140248006733216: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006733216: core_fifo_inputs_t;
        signal outputs_full_140248006733216: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006733272: core_fifo_inputs_t;
        signal fifo_full_140248006733272: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006733272: core_fifo_inputs_t;
        signal outputs_full_140248006733272: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006733328: core_fifo_inputs_t;
        signal fifo_full_140248006733328: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006733328: core_fifo_inputs_t;
        signal outputs_full_140248006733328: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006733384: core_fifo_inputs_t;
        signal fifo_full_140248006733384: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006733384: core_fifo_inputs_t;
        signal outputs_full_140248006733384: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006733440: core_fifo_inputs_t;
        signal fifo_full_140248006733440: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006733440: core_fifo_inputs_t;
        signal outputs_full_140248006733440: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006733496: core_fifo_inputs_t;
        signal fifo_full_140248006733496: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006733496: core_fifo_inputs_t;
        signal outputs_full_140248006733496: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006733552: core_fifo_inputs_t;
        signal fifo_full_140248006733552: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006733552: core_fifo_inputs_t;
        signal outputs_full_140248006733552: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006733608: core_fifo_inputs_t;
        signal fifo_full_140248006733608: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006733608: core_fifo_inputs_t;
        signal outputs_full_140248006733608: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006733664: core_fifo_inputs_t;
        signal fifo_full_140248006733664: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006733664: core_fifo_inputs_t;
        signal outputs_full_140248006733664: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006733720: core_fifo_inputs_t;
        signal fifo_full_140248006733720: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006733720: core_fifo_inputs_t;
        signal outputs_full_140248006733720: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006733776: core_fifo_inputs_t;
        signal fifo_full_140248006733776: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006733776: core_fifo_inputs_t;
        signal outputs_full_140248006733776: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006750280: core_fifo_inputs_t;
        signal fifo_full_140248006750280: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006750280: core_fifo_inputs_t;
        signal outputs_full_140248006750280: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006750336: core_fifo_inputs_t;
        signal fifo_full_140248006750336: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006750336: core_fifo_inputs_t;
        signal outputs_full_140248006750336: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006750392: core_fifo_inputs_t;
        signal fifo_full_140248006750392: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006750392: core_fifo_inputs_t;
        signal outputs_full_140248006750392: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006750448: core_fifo_inputs_t;
        signal fifo_full_140248006750448: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006750448: core_fifo_inputs_t;
        signal outputs_full_140248006750448: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006750504: core_fifo_inputs_t;
        signal fifo_full_140248006750504: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006750504: core_fifo_inputs_t;
        signal outputs_full_140248006750504: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006750560: core_fifo_inputs_t;
        signal fifo_full_140248006750560: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006750560: core_fifo_inputs_t;
        signal outputs_full_140248006750560: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006750616: core_fifo_inputs_t;
        signal fifo_full_140248006750616: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006750616: core_fifo_inputs_t;
        signal outputs_full_140248006750616: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006750672: core_fifo_inputs_t;
        signal fifo_full_140248006750672: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006750672: core_fifo_inputs_t;
        signal outputs_full_140248006750672: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006750728: core_fifo_inputs_t;
        signal fifo_full_140248006750728: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006750728: core_fifo_inputs_t;
        signal outputs_full_140248006750728: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006750784: core_fifo_inputs_t;
        signal fifo_full_140248006750784: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006750784: core_fifo_inputs_t;
        signal outputs_full_140248006750784: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006750840: core_fifo_inputs_t;
        signal fifo_full_140248006750840: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006750840: core_fifo_inputs_t;
        signal outputs_full_140248006750840: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006750896: core_fifo_inputs_t;
        signal fifo_full_140248006750896: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006750896: core_fifo_inputs_t;
        signal outputs_full_140248006750896: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006750952: core_fifo_inputs_t;
        signal fifo_full_140248006750952: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006750952: core_fifo_inputs_t;
        signal outputs_full_140248006750952: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006751008: core_fifo_inputs_t;
        signal fifo_full_140248006751008: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006751008: core_fifo_inputs_t;
        signal outputs_full_140248006751008: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006751064: core_fifo_inputs_t;
        signal fifo_full_140248006751064: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006751064: core_fifo_inputs_t;
        signal outputs_full_140248006751064: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006751120: core_fifo_inputs_t;
        signal fifo_full_140248006751120: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006751120: core_fifo_inputs_t;
        signal outputs_full_140248006751120: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006751176: core_fifo_inputs_t;
        signal fifo_full_140248006751176: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006751176: core_fifo_inputs_t;
        signal outputs_full_140248006751176: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006751232: core_fifo_inputs_t;
        signal fifo_full_140248006751232: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006751232: core_fifo_inputs_t;
        signal outputs_full_140248006751232: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006751288: core_fifo_inputs_t;
        signal fifo_full_140248006751288: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006751288: core_fifo_inputs_t;
        signal outputs_full_140248006751288: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006751344: core_fifo_inputs_t;
        signal fifo_full_140248006751344: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006751344: core_fifo_inputs_t;
        signal outputs_full_140248006751344: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006751400: core_fifo_inputs_t;
        signal fifo_full_140248006751400: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006751400: core_fifo_inputs_t;
        signal outputs_full_140248006751400: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006751456: core_fifo_inputs_t;
        signal fifo_full_140248006751456: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006751456: core_fifo_inputs_t;
        signal outputs_full_140248006751456: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006751512: core_fifo_inputs_t;
        signal fifo_full_140248006751512: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006751512: core_fifo_inputs_t;
        signal outputs_full_140248006751512: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006751568: core_fifo_inputs_t;
        signal fifo_full_140248006751568: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006751568: core_fifo_inputs_t;
        signal outputs_full_140248006751568: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006751624: core_fifo_inputs_t;
        signal fifo_full_140248006751624: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006751624: core_fifo_inputs_t;
        signal outputs_full_140248006751624: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006751680: core_fifo_inputs_t;
        signal fifo_full_140248006751680: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006751680: core_fifo_inputs_t;
        signal outputs_full_140248006751680: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006751736: core_fifo_inputs_t;
        signal fifo_full_140248006751736: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006751736: core_fifo_inputs_t;
        signal outputs_full_140248006751736: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006751792: core_fifo_inputs_t;
        signal fifo_full_140248006751792: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006751792: core_fifo_inputs_t;
        signal outputs_full_140248006751792: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006751848: core_fifo_inputs_t;
        signal fifo_full_140248006751848: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006751848: core_fifo_inputs_t;
        signal outputs_full_140248006751848: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006751904: core_fifo_inputs_t;
        signal fifo_full_140248006751904: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006751904: core_fifo_inputs_t;
        signal outputs_full_140248006751904: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006751960: core_fifo_inputs_t;
        signal fifo_full_140248006751960: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006751960: core_fifo_inputs_t;
        signal outputs_full_140248006751960: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006752016: core_fifo_inputs_t;
        signal fifo_full_140248006752016: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006752016: core_fifo_inputs_t;
        signal outputs_full_140248006752016: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006752072: core_fifo_inputs_t;
        signal fifo_full_140248006752072: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006752072: core_fifo_inputs_t;
        signal outputs_full_140248006752072: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006752128: core_fifo_inputs_t;
        signal fifo_full_140248006752128: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006752128: core_fifo_inputs_t;
        signal outputs_full_140248006752128: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006752184: core_fifo_inputs_t;
        signal fifo_full_140248006752184: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006752184: core_fifo_inputs_t;
        signal outputs_full_140248006752184: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006752240: core_fifo_inputs_t;
        signal fifo_full_140248006752240: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006752240: core_fifo_inputs_t;
        signal outputs_full_140248006752240: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006752296: core_fifo_inputs_t;
        signal fifo_full_140248006752296: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006752296: core_fifo_inputs_t;
        signal outputs_full_140248006752296: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006752352: core_fifo_inputs_t;
        signal fifo_full_140248006752352: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006752352: core_fifo_inputs_t;
        signal outputs_full_140248006752352: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_140248006752408: core_fifo_inputs_t;
        signal fifo_full_140248006752408: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_140248006752408: core_fifo_inputs_t;
        signal outputs_full_140248006752408: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        

begin

        outputs(0) <= outputs_140248006752408(0);
        outputs_full_140248006752408(0) <= outputs_full(0);
        
        outputs(1) <= outputs_140248006679688(1);
        outputs_full_140248006679688(1) <= outputs_full(1);
        
        fifo_inputs_140248006752408(0) <= fifo_inputs(0);
        fifo_full(0) <= fifo_full_140248006752408(0);
                
        fifo_inputs_140248006679688(1) <= fifo_inputs(1);
        fifo_full(1) <= fifo_full_140248006679688(1);
    
        fifo_inputs_140248006679632(1) <= outputs_140248006679688(0);
        outputs_full_140248006679688(0) <= fifo_full_140248006679632(1);
        
        fifo_inputs_140248006679856(1) <= outputs_140248006679632(0);
        outputs_full_140248006679632(0) <= fifo_full_140248006679856(1);
        
        fifo_inputs_140248006679688(0) <= outputs_140248006679632(1);
        outputs_full_140248006679632(1) <= fifo_full_140248006679688(0);
        
        fifo_inputs_140248006679912(1) <= outputs_140248006679856(0);
        outputs_full_140248006679856(0) <= fifo_full_140248006679912(1);
        
        fifo_inputs_140248006679632(0) <= outputs_140248006679856(1);
        outputs_full_140248006679856(1) <= fifo_full_140248006679632(0);
        
        fifo_inputs_140248006679968(1) <= outputs_140248006679912(0);
        outputs_full_140248006679912(0) <= fifo_full_140248006679968(1);
        
        fifo_inputs_140248006679856(0) <= outputs_140248006679912(1);
        outputs_full_140248006679912(1) <= fifo_full_140248006679856(0);
        
        fifo_inputs_140248006679800(1) <= outputs_140248006679968(0);
        outputs_full_140248006679968(0) <= fifo_full_140248006679800(1);
        
        fifo_inputs_140248006679912(0) <= outputs_140248006679968(1);
        outputs_full_140248006679968(1) <= fifo_full_140248006679912(0);
        
        fifo_inputs_140248006680024(1) <= outputs_140248006679800(0);
        outputs_full_140248006679800(0) <= fifo_full_140248006680024(1);
        
        fifo_inputs_140248006679968(0) <= outputs_140248006679800(1);
        outputs_full_140248006679800(1) <= fifo_full_140248006679968(0);
        
        fifo_inputs_140248006680080(1) <= outputs_140248006680024(0);
        outputs_full_140248006680024(0) <= fifo_full_140248006680080(1);
        
        fifo_inputs_140248006679800(0) <= outputs_140248006680024(1);
        outputs_full_140248006680024(1) <= fifo_full_140248006679800(0);
        
        fifo_inputs_140248006680136(1) <= outputs_140248006680080(0);
        outputs_full_140248006680080(0) <= fifo_full_140248006680136(1);
        
        fifo_inputs_140248006680024(0) <= outputs_140248006680080(1);
        outputs_full_140248006680080(1) <= fifo_full_140248006680024(0);
        
        fifo_inputs_140248006680192(1) <= outputs_140248006680136(0);
        outputs_full_140248006680136(0) <= fifo_full_140248006680192(1);
        
        fifo_inputs_140248006680080(0) <= outputs_140248006680136(1);
        outputs_full_140248006680136(1) <= fifo_full_140248006680080(0);
        
        fifo_inputs_140248006679744(1) <= outputs_140248006680192(0);
        outputs_full_140248006680192(0) <= fifo_full_140248006679744(1);
        
        fifo_inputs_140248006680136(0) <= outputs_140248006680192(1);
        outputs_full_140248006680192(1) <= fifo_full_140248006680136(0);
        
        fifo_inputs_140248006680248(1) <= outputs_140248006679744(0);
        outputs_full_140248006679744(0) <= fifo_full_140248006680248(1);
        
        fifo_inputs_140248006680192(0) <= outputs_140248006679744(1);
        outputs_full_140248006679744(1) <= fifo_full_140248006680192(0);
        
        fifo_inputs_140248006680304(1) <= outputs_140248006680248(0);
        outputs_full_140248006680248(0) <= fifo_full_140248006680304(1);
        
        fifo_inputs_140248006679744(0) <= outputs_140248006680248(1);
        outputs_full_140248006680248(1) <= fifo_full_140248006679744(0);
        
        fifo_inputs_140248006680360(1) <= outputs_140248006680304(0);
        outputs_full_140248006680304(0) <= fifo_full_140248006680360(1);
        
        fifo_inputs_140248006680248(0) <= outputs_140248006680304(1);
        outputs_full_140248006680304(1) <= fifo_full_140248006680248(0);
        
        fifo_inputs_140248006680416(1) <= outputs_140248006680360(0);
        outputs_full_140248006680360(0) <= fifo_full_140248006680416(1);
        
        fifo_inputs_140248006680304(0) <= outputs_140248006680360(1);
        outputs_full_140248006680360(1) <= fifo_full_140248006680304(0);
        
        fifo_inputs_140248006680472(1) <= outputs_140248006680416(0);
        outputs_full_140248006680416(0) <= fifo_full_140248006680472(1);
        
        fifo_inputs_140248006680360(0) <= outputs_140248006680416(1);
        outputs_full_140248006680416(1) <= fifo_full_140248006680360(0);
        
        fifo_inputs_140248006680528(1) <= outputs_140248006680472(0);
        outputs_full_140248006680472(0) <= fifo_full_140248006680528(1);
        
        fifo_inputs_140248006680416(0) <= outputs_140248006680472(1);
        outputs_full_140248006680472(1) <= fifo_full_140248006680416(0);
        
        fifo_inputs_140248006729800(1) <= outputs_140248006680528(0);
        outputs_full_140248006680528(0) <= fifo_full_140248006729800(1);
        
        fifo_inputs_140248006680472(0) <= outputs_140248006680528(1);
        outputs_full_140248006680528(1) <= fifo_full_140248006680472(0);
        
        fifo_inputs_140248006729856(1) <= outputs_140248006729800(0);
        outputs_full_140248006729800(0) <= fifo_full_140248006729856(1);
        
        fifo_inputs_140248006680528(0) <= outputs_140248006729800(1);
        outputs_full_140248006729800(1) <= fifo_full_140248006680528(0);
        
        fifo_inputs_140248006729912(1) <= outputs_140248006729856(0);
        outputs_full_140248006729856(0) <= fifo_full_140248006729912(1);
        
        fifo_inputs_140248006729800(0) <= outputs_140248006729856(1);
        outputs_full_140248006729856(1) <= fifo_full_140248006729800(0);
        
        fifo_inputs_140248006729968(1) <= outputs_140248006729912(0);
        outputs_full_140248006729912(0) <= fifo_full_140248006729968(1);
        
        fifo_inputs_140248006729856(0) <= outputs_140248006729912(1);
        outputs_full_140248006729912(1) <= fifo_full_140248006729856(0);
        
        fifo_inputs_140248006730024(1) <= outputs_140248006729968(0);
        outputs_full_140248006729968(0) <= fifo_full_140248006730024(1);
        
        fifo_inputs_140248006729912(0) <= outputs_140248006729968(1);
        outputs_full_140248006729968(1) <= fifo_full_140248006729912(0);
        
        fifo_inputs_140248006730080(1) <= outputs_140248006730024(0);
        outputs_full_140248006730024(0) <= fifo_full_140248006730080(1);
        
        fifo_inputs_140248006729968(0) <= outputs_140248006730024(1);
        outputs_full_140248006730024(1) <= fifo_full_140248006729968(0);
        
        fifo_inputs_140248006730136(1) <= outputs_140248006730080(0);
        outputs_full_140248006730080(0) <= fifo_full_140248006730136(1);
        
        fifo_inputs_140248006730024(0) <= outputs_140248006730080(1);
        outputs_full_140248006730080(1) <= fifo_full_140248006730024(0);
        
        fifo_inputs_140248006730192(1) <= outputs_140248006730136(0);
        outputs_full_140248006730136(0) <= fifo_full_140248006730192(1);
        
        fifo_inputs_140248006730080(0) <= outputs_140248006730136(1);
        outputs_full_140248006730136(1) <= fifo_full_140248006730080(0);
        
        fifo_inputs_140248006730248(1) <= outputs_140248006730192(0);
        outputs_full_140248006730192(0) <= fifo_full_140248006730248(1);
        
        fifo_inputs_140248006730136(0) <= outputs_140248006730192(1);
        outputs_full_140248006730192(1) <= fifo_full_140248006730136(0);
        
        fifo_inputs_140248006730304(1) <= outputs_140248006730248(0);
        outputs_full_140248006730248(0) <= fifo_full_140248006730304(1);
        
        fifo_inputs_140248006730192(0) <= outputs_140248006730248(1);
        outputs_full_140248006730248(1) <= fifo_full_140248006730192(0);
        
        fifo_inputs_140248006730360(1) <= outputs_140248006730304(0);
        outputs_full_140248006730304(0) <= fifo_full_140248006730360(1);
        
        fifo_inputs_140248006730248(0) <= outputs_140248006730304(1);
        outputs_full_140248006730304(1) <= fifo_full_140248006730248(0);
        
        fifo_inputs_140248006730416(1) <= outputs_140248006730360(0);
        outputs_full_140248006730360(0) <= fifo_full_140248006730416(1);
        
        fifo_inputs_140248006730304(0) <= outputs_140248006730360(1);
        outputs_full_140248006730360(1) <= fifo_full_140248006730304(0);
        
        fifo_inputs_140248006730472(1) <= outputs_140248006730416(0);
        outputs_full_140248006730416(0) <= fifo_full_140248006730472(1);
        
        fifo_inputs_140248006730360(0) <= outputs_140248006730416(1);
        outputs_full_140248006730416(1) <= fifo_full_140248006730360(0);
        
        fifo_inputs_140248006730528(1) <= outputs_140248006730472(0);
        outputs_full_140248006730472(0) <= fifo_full_140248006730528(1);
        
        fifo_inputs_140248006730416(0) <= outputs_140248006730472(1);
        outputs_full_140248006730472(1) <= fifo_full_140248006730416(0);
        
        fifo_inputs_140248006730584(1) <= outputs_140248006730528(0);
        outputs_full_140248006730528(0) <= fifo_full_140248006730584(1);
        
        fifo_inputs_140248006730472(0) <= outputs_140248006730528(1);
        outputs_full_140248006730528(1) <= fifo_full_140248006730472(0);
        
        fifo_inputs_140248006730640(1) <= outputs_140248006730584(0);
        outputs_full_140248006730584(0) <= fifo_full_140248006730640(1);
        
        fifo_inputs_140248006730528(0) <= outputs_140248006730584(1);
        outputs_full_140248006730584(1) <= fifo_full_140248006730528(0);
        
        fifo_inputs_140248006730696(1) <= outputs_140248006730640(0);
        outputs_full_140248006730640(0) <= fifo_full_140248006730696(1);
        
        fifo_inputs_140248006730584(0) <= outputs_140248006730640(1);
        outputs_full_140248006730640(1) <= fifo_full_140248006730584(0);
        
        fifo_inputs_140248006730752(1) <= outputs_140248006730696(0);
        outputs_full_140248006730696(0) <= fifo_full_140248006730752(1);
        
        fifo_inputs_140248006730640(0) <= outputs_140248006730696(1);
        outputs_full_140248006730696(1) <= fifo_full_140248006730640(0);
        
        fifo_inputs_140248006730808(1) <= outputs_140248006730752(0);
        outputs_full_140248006730752(0) <= fifo_full_140248006730808(1);
        
        fifo_inputs_140248006730696(0) <= outputs_140248006730752(1);
        outputs_full_140248006730752(1) <= fifo_full_140248006730696(0);
        
        fifo_inputs_140248006730864(1) <= outputs_140248006730808(0);
        outputs_full_140248006730808(0) <= fifo_full_140248006730864(1);
        
        fifo_inputs_140248006730752(0) <= outputs_140248006730808(1);
        outputs_full_140248006730808(1) <= fifo_full_140248006730752(0);
        
        fifo_inputs_140248006730920(1) <= outputs_140248006730864(0);
        outputs_full_140248006730864(0) <= fifo_full_140248006730920(1);
        
        fifo_inputs_140248006730808(0) <= outputs_140248006730864(1);
        outputs_full_140248006730864(1) <= fifo_full_140248006730808(0);
        
        fifo_inputs_140248006730976(1) <= outputs_140248006730920(0);
        outputs_full_140248006730920(0) <= fifo_full_140248006730976(1);
        
        fifo_inputs_140248006730864(0) <= outputs_140248006730920(1);
        outputs_full_140248006730920(1) <= fifo_full_140248006730864(0);
        
        fifo_inputs_140248006731032(1) <= outputs_140248006730976(0);
        outputs_full_140248006730976(0) <= fifo_full_140248006731032(1);
        
        fifo_inputs_140248006730920(0) <= outputs_140248006730976(1);
        outputs_full_140248006730976(1) <= fifo_full_140248006730920(0);
        
        fifo_inputs_140248006731088(1) <= outputs_140248006731032(0);
        outputs_full_140248006731032(0) <= fifo_full_140248006731088(1);
        
        fifo_inputs_140248006730976(0) <= outputs_140248006731032(1);
        outputs_full_140248006731032(1) <= fifo_full_140248006730976(0);
        
        fifo_inputs_140248006731144(1) <= outputs_140248006731088(0);
        outputs_full_140248006731088(0) <= fifo_full_140248006731144(1);
        
        fifo_inputs_140248006731032(0) <= outputs_140248006731088(1);
        outputs_full_140248006731088(1) <= fifo_full_140248006731032(0);
        
        fifo_inputs_140248006731200(1) <= outputs_140248006731144(0);
        outputs_full_140248006731144(0) <= fifo_full_140248006731200(1);
        
        fifo_inputs_140248006731088(0) <= outputs_140248006731144(1);
        outputs_full_140248006731144(1) <= fifo_full_140248006731088(0);
        
        fifo_inputs_140248006731256(1) <= outputs_140248006731200(0);
        outputs_full_140248006731200(0) <= fifo_full_140248006731256(1);
        
        fifo_inputs_140248006731144(0) <= outputs_140248006731200(1);
        outputs_full_140248006731200(1) <= fifo_full_140248006731144(0);
        
        fifo_inputs_140248006731312(1) <= outputs_140248006731256(0);
        outputs_full_140248006731256(0) <= fifo_full_140248006731312(1);
        
        fifo_inputs_140248006731200(0) <= outputs_140248006731256(1);
        outputs_full_140248006731256(1) <= fifo_full_140248006731200(0);
        
        fifo_inputs_140248006731368(1) <= outputs_140248006731312(0);
        outputs_full_140248006731312(0) <= fifo_full_140248006731368(1);
        
        fifo_inputs_140248006731256(0) <= outputs_140248006731312(1);
        outputs_full_140248006731312(1) <= fifo_full_140248006731256(0);
        
        fifo_inputs_140248006731424(1) <= outputs_140248006731368(0);
        outputs_full_140248006731368(0) <= fifo_full_140248006731424(1);
        
        fifo_inputs_140248006731312(0) <= outputs_140248006731368(1);
        outputs_full_140248006731368(1) <= fifo_full_140248006731312(0);
        
        fifo_inputs_140248006731480(1) <= outputs_140248006731424(0);
        outputs_full_140248006731424(0) <= fifo_full_140248006731480(1);
        
        fifo_inputs_140248006731368(0) <= outputs_140248006731424(1);
        outputs_full_140248006731424(1) <= fifo_full_140248006731368(0);
        
        fifo_inputs_140248006731536(1) <= outputs_140248006731480(0);
        outputs_full_140248006731480(0) <= fifo_full_140248006731536(1);
        
        fifo_inputs_140248006731424(0) <= outputs_140248006731480(1);
        outputs_full_140248006731480(1) <= fifo_full_140248006731424(0);
        
        fifo_inputs_140248006731592(1) <= outputs_140248006731536(0);
        outputs_full_140248006731536(0) <= fifo_full_140248006731592(1);
        
        fifo_inputs_140248006731480(0) <= outputs_140248006731536(1);
        outputs_full_140248006731536(1) <= fifo_full_140248006731480(0);
        
        fifo_inputs_140248006731648(1) <= outputs_140248006731592(0);
        outputs_full_140248006731592(0) <= fifo_full_140248006731648(1);
        
        fifo_inputs_140248006731536(0) <= outputs_140248006731592(1);
        outputs_full_140248006731592(1) <= fifo_full_140248006731536(0);
        
        fifo_inputs_140248006731704(1) <= outputs_140248006731648(0);
        outputs_full_140248006731648(0) <= fifo_full_140248006731704(1);
        
        fifo_inputs_140248006731592(0) <= outputs_140248006731648(1);
        outputs_full_140248006731648(1) <= fifo_full_140248006731592(0);
        
        fifo_inputs_140248006731760(1) <= outputs_140248006731704(0);
        outputs_full_140248006731704(0) <= fifo_full_140248006731760(1);
        
        fifo_inputs_140248006731648(0) <= outputs_140248006731704(1);
        outputs_full_140248006731704(1) <= fifo_full_140248006731648(0);
        
        fifo_inputs_140248006731816(1) <= outputs_140248006731760(0);
        outputs_full_140248006731760(0) <= fifo_full_140248006731816(1);
        
        fifo_inputs_140248006731704(0) <= outputs_140248006731760(1);
        outputs_full_140248006731760(1) <= fifo_full_140248006731704(0);
        
        fifo_inputs_140248006731872(1) <= outputs_140248006731816(0);
        outputs_full_140248006731816(0) <= fifo_full_140248006731872(1);
        
        fifo_inputs_140248006731760(0) <= outputs_140248006731816(1);
        outputs_full_140248006731816(1) <= fifo_full_140248006731760(0);
        
        fifo_inputs_140248006731928(1) <= outputs_140248006731872(0);
        outputs_full_140248006731872(0) <= fifo_full_140248006731928(1);
        
        fifo_inputs_140248006731816(0) <= outputs_140248006731872(1);
        outputs_full_140248006731872(1) <= fifo_full_140248006731816(0);
        
        fifo_inputs_140248006731984(1) <= outputs_140248006731928(0);
        outputs_full_140248006731928(0) <= fifo_full_140248006731984(1);
        
        fifo_inputs_140248006731872(0) <= outputs_140248006731928(1);
        outputs_full_140248006731928(1) <= fifo_full_140248006731872(0);
        
        fifo_inputs_140248006732040(1) <= outputs_140248006731984(0);
        outputs_full_140248006731984(0) <= fifo_full_140248006732040(1);
        
        fifo_inputs_140248006731928(0) <= outputs_140248006731984(1);
        outputs_full_140248006731984(1) <= fifo_full_140248006731928(0);
        
        fifo_inputs_140248006732096(1) <= outputs_140248006732040(0);
        outputs_full_140248006732040(0) <= fifo_full_140248006732096(1);
        
        fifo_inputs_140248006731984(0) <= outputs_140248006732040(1);
        outputs_full_140248006732040(1) <= fifo_full_140248006731984(0);
        
        fifo_inputs_140248006732152(1) <= outputs_140248006732096(0);
        outputs_full_140248006732096(0) <= fifo_full_140248006732152(1);
        
        fifo_inputs_140248006732040(0) <= outputs_140248006732096(1);
        outputs_full_140248006732096(1) <= fifo_full_140248006732040(0);
        
        fifo_inputs_140248006732208(1) <= outputs_140248006732152(0);
        outputs_full_140248006732152(0) <= fifo_full_140248006732208(1);
        
        fifo_inputs_140248006732096(0) <= outputs_140248006732152(1);
        outputs_full_140248006732152(1) <= fifo_full_140248006732096(0);
        
        fifo_inputs_140248006732264(1) <= outputs_140248006732208(0);
        outputs_full_140248006732208(0) <= fifo_full_140248006732264(1);
        
        fifo_inputs_140248006732152(0) <= outputs_140248006732208(1);
        outputs_full_140248006732208(1) <= fifo_full_140248006732152(0);
        
        fifo_inputs_140248006732320(1) <= outputs_140248006732264(0);
        outputs_full_140248006732264(0) <= fifo_full_140248006732320(1);
        
        fifo_inputs_140248006732208(0) <= outputs_140248006732264(1);
        outputs_full_140248006732264(1) <= fifo_full_140248006732208(0);
        
        fifo_inputs_140248006732376(1) <= outputs_140248006732320(0);
        outputs_full_140248006732320(0) <= fifo_full_140248006732376(1);
        
        fifo_inputs_140248006732264(0) <= outputs_140248006732320(1);
        outputs_full_140248006732320(1) <= fifo_full_140248006732264(0);
        
        fifo_inputs_140248006732432(1) <= outputs_140248006732376(0);
        outputs_full_140248006732376(0) <= fifo_full_140248006732432(1);
        
        fifo_inputs_140248006732320(0) <= outputs_140248006732376(1);
        outputs_full_140248006732376(1) <= fifo_full_140248006732320(0);
        
        fifo_inputs_140248006732488(1) <= outputs_140248006732432(0);
        outputs_full_140248006732432(0) <= fifo_full_140248006732488(1);
        
        fifo_inputs_140248006732376(0) <= outputs_140248006732432(1);
        outputs_full_140248006732432(1) <= fifo_full_140248006732376(0);
        
        fifo_inputs_140248006732544(1) <= outputs_140248006732488(0);
        outputs_full_140248006732488(0) <= fifo_full_140248006732544(1);
        
        fifo_inputs_140248006732432(0) <= outputs_140248006732488(1);
        outputs_full_140248006732488(1) <= fifo_full_140248006732432(0);
        
        fifo_inputs_140248006732600(1) <= outputs_140248006732544(0);
        outputs_full_140248006732544(0) <= fifo_full_140248006732600(1);
        
        fifo_inputs_140248006732488(0) <= outputs_140248006732544(1);
        outputs_full_140248006732544(1) <= fifo_full_140248006732488(0);
        
        fifo_inputs_140248006732656(1) <= outputs_140248006732600(0);
        outputs_full_140248006732600(0) <= fifo_full_140248006732656(1);
        
        fifo_inputs_140248006732544(0) <= outputs_140248006732600(1);
        outputs_full_140248006732600(1) <= fifo_full_140248006732544(0);
        
        fifo_inputs_140248006732712(1) <= outputs_140248006732656(0);
        outputs_full_140248006732656(0) <= fifo_full_140248006732712(1);
        
        fifo_inputs_140248006732600(0) <= outputs_140248006732656(1);
        outputs_full_140248006732656(1) <= fifo_full_140248006732600(0);
        
        fifo_inputs_140248006732768(1) <= outputs_140248006732712(0);
        outputs_full_140248006732712(0) <= fifo_full_140248006732768(1);
        
        fifo_inputs_140248006732656(0) <= outputs_140248006732712(1);
        outputs_full_140248006732712(1) <= fifo_full_140248006732656(0);
        
        fifo_inputs_140248006732824(1) <= outputs_140248006732768(0);
        outputs_full_140248006732768(0) <= fifo_full_140248006732824(1);
        
        fifo_inputs_140248006732712(0) <= outputs_140248006732768(1);
        outputs_full_140248006732768(1) <= fifo_full_140248006732712(0);
        
        fifo_inputs_140248006732880(1) <= outputs_140248006732824(0);
        outputs_full_140248006732824(0) <= fifo_full_140248006732880(1);
        
        fifo_inputs_140248006732768(0) <= outputs_140248006732824(1);
        outputs_full_140248006732824(1) <= fifo_full_140248006732768(0);
        
        fifo_inputs_140248006732936(1) <= outputs_140248006732880(0);
        outputs_full_140248006732880(0) <= fifo_full_140248006732936(1);
        
        fifo_inputs_140248006732824(0) <= outputs_140248006732880(1);
        outputs_full_140248006732880(1) <= fifo_full_140248006732824(0);
        
        fifo_inputs_140248006732992(1) <= outputs_140248006732936(0);
        outputs_full_140248006732936(0) <= fifo_full_140248006732992(1);
        
        fifo_inputs_140248006732880(0) <= outputs_140248006732936(1);
        outputs_full_140248006732936(1) <= fifo_full_140248006732880(0);
        
        fifo_inputs_140248006733048(1) <= outputs_140248006732992(0);
        outputs_full_140248006732992(0) <= fifo_full_140248006733048(1);
        
        fifo_inputs_140248006732936(0) <= outputs_140248006732992(1);
        outputs_full_140248006732992(1) <= fifo_full_140248006732936(0);
        
        fifo_inputs_140248006733104(1) <= outputs_140248006733048(0);
        outputs_full_140248006733048(0) <= fifo_full_140248006733104(1);
        
        fifo_inputs_140248006732992(0) <= outputs_140248006733048(1);
        outputs_full_140248006733048(1) <= fifo_full_140248006732992(0);
        
        fifo_inputs_140248006733160(1) <= outputs_140248006733104(0);
        outputs_full_140248006733104(0) <= fifo_full_140248006733160(1);
        
        fifo_inputs_140248006733048(0) <= outputs_140248006733104(1);
        outputs_full_140248006733104(1) <= fifo_full_140248006733048(0);
        
        fifo_inputs_140248006733216(1) <= outputs_140248006733160(0);
        outputs_full_140248006733160(0) <= fifo_full_140248006733216(1);
        
        fifo_inputs_140248006733104(0) <= outputs_140248006733160(1);
        outputs_full_140248006733160(1) <= fifo_full_140248006733104(0);
        
        fifo_inputs_140248006733272(1) <= outputs_140248006733216(0);
        outputs_full_140248006733216(0) <= fifo_full_140248006733272(1);
        
        fifo_inputs_140248006733160(0) <= outputs_140248006733216(1);
        outputs_full_140248006733216(1) <= fifo_full_140248006733160(0);
        
        fifo_inputs_140248006733328(1) <= outputs_140248006733272(0);
        outputs_full_140248006733272(0) <= fifo_full_140248006733328(1);
        
        fifo_inputs_140248006733216(0) <= outputs_140248006733272(1);
        outputs_full_140248006733272(1) <= fifo_full_140248006733216(0);
        
        fifo_inputs_140248006733384(1) <= outputs_140248006733328(0);
        outputs_full_140248006733328(0) <= fifo_full_140248006733384(1);
        
        fifo_inputs_140248006733272(0) <= outputs_140248006733328(1);
        outputs_full_140248006733328(1) <= fifo_full_140248006733272(0);
        
        fifo_inputs_140248006733440(1) <= outputs_140248006733384(0);
        outputs_full_140248006733384(0) <= fifo_full_140248006733440(1);
        
        fifo_inputs_140248006733328(0) <= outputs_140248006733384(1);
        outputs_full_140248006733384(1) <= fifo_full_140248006733328(0);
        
        fifo_inputs_140248006733496(1) <= outputs_140248006733440(0);
        outputs_full_140248006733440(0) <= fifo_full_140248006733496(1);
        
        fifo_inputs_140248006733384(0) <= outputs_140248006733440(1);
        outputs_full_140248006733440(1) <= fifo_full_140248006733384(0);
        
        fifo_inputs_140248006733552(1) <= outputs_140248006733496(0);
        outputs_full_140248006733496(0) <= fifo_full_140248006733552(1);
        
        fifo_inputs_140248006733440(0) <= outputs_140248006733496(1);
        outputs_full_140248006733496(1) <= fifo_full_140248006733440(0);
        
        fifo_inputs_140248006733608(1) <= outputs_140248006733552(0);
        outputs_full_140248006733552(0) <= fifo_full_140248006733608(1);
        
        fifo_inputs_140248006733496(0) <= outputs_140248006733552(1);
        outputs_full_140248006733552(1) <= fifo_full_140248006733496(0);
        
        fifo_inputs_140248006733664(1) <= outputs_140248006733608(0);
        outputs_full_140248006733608(0) <= fifo_full_140248006733664(1);
        
        fifo_inputs_140248006733552(0) <= outputs_140248006733608(1);
        outputs_full_140248006733608(1) <= fifo_full_140248006733552(0);
        
        fifo_inputs_140248006733720(1) <= outputs_140248006733664(0);
        outputs_full_140248006733664(0) <= fifo_full_140248006733720(1);
        
        fifo_inputs_140248006733608(0) <= outputs_140248006733664(1);
        outputs_full_140248006733664(1) <= fifo_full_140248006733608(0);
        
        fifo_inputs_140248006733776(1) <= outputs_140248006733720(0);
        outputs_full_140248006733720(0) <= fifo_full_140248006733776(1);
        
        fifo_inputs_140248006733664(0) <= outputs_140248006733720(1);
        outputs_full_140248006733720(1) <= fifo_full_140248006733664(0);
        
        fifo_inputs_140248006750280(1) <= outputs_140248006733776(0);
        outputs_full_140248006733776(0) <= fifo_full_140248006750280(1);
        
        fifo_inputs_140248006733720(0) <= outputs_140248006733776(1);
        outputs_full_140248006733776(1) <= fifo_full_140248006733720(0);
        
        fifo_inputs_140248006750336(1) <= outputs_140248006750280(0);
        outputs_full_140248006750280(0) <= fifo_full_140248006750336(1);
        
        fifo_inputs_140248006733776(0) <= outputs_140248006750280(1);
        outputs_full_140248006750280(1) <= fifo_full_140248006733776(0);
        
        fifo_inputs_140248006750392(1) <= outputs_140248006750336(0);
        outputs_full_140248006750336(0) <= fifo_full_140248006750392(1);
        
        fifo_inputs_140248006750280(0) <= outputs_140248006750336(1);
        outputs_full_140248006750336(1) <= fifo_full_140248006750280(0);
        
        fifo_inputs_140248006750448(1) <= outputs_140248006750392(0);
        outputs_full_140248006750392(0) <= fifo_full_140248006750448(1);
        
        fifo_inputs_140248006750336(0) <= outputs_140248006750392(1);
        outputs_full_140248006750392(1) <= fifo_full_140248006750336(0);
        
        fifo_inputs_140248006750504(1) <= outputs_140248006750448(0);
        outputs_full_140248006750448(0) <= fifo_full_140248006750504(1);
        
        fifo_inputs_140248006750392(0) <= outputs_140248006750448(1);
        outputs_full_140248006750448(1) <= fifo_full_140248006750392(0);
        
        fifo_inputs_140248006750560(1) <= outputs_140248006750504(0);
        outputs_full_140248006750504(0) <= fifo_full_140248006750560(1);
        
        fifo_inputs_140248006750448(0) <= outputs_140248006750504(1);
        outputs_full_140248006750504(1) <= fifo_full_140248006750448(0);
        
        fifo_inputs_140248006750616(1) <= outputs_140248006750560(0);
        outputs_full_140248006750560(0) <= fifo_full_140248006750616(1);
        
        fifo_inputs_140248006750504(0) <= outputs_140248006750560(1);
        outputs_full_140248006750560(1) <= fifo_full_140248006750504(0);
        
        fifo_inputs_140248006750672(1) <= outputs_140248006750616(0);
        outputs_full_140248006750616(0) <= fifo_full_140248006750672(1);
        
        fifo_inputs_140248006750560(0) <= outputs_140248006750616(1);
        outputs_full_140248006750616(1) <= fifo_full_140248006750560(0);
        
        fifo_inputs_140248006750728(1) <= outputs_140248006750672(0);
        outputs_full_140248006750672(0) <= fifo_full_140248006750728(1);
        
        fifo_inputs_140248006750616(0) <= outputs_140248006750672(1);
        outputs_full_140248006750672(1) <= fifo_full_140248006750616(0);
        
        fifo_inputs_140248006750784(1) <= outputs_140248006750728(0);
        outputs_full_140248006750728(0) <= fifo_full_140248006750784(1);
        
        fifo_inputs_140248006750672(0) <= outputs_140248006750728(1);
        outputs_full_140248006750728(1) <= fifo_full_140248006750672(0);
        
        fifo_inputs_140248006750840(1) <= outputs_140248006750784(0);
        outputs_full_140248006750784(0) <= fifo_full_140248006750840(1);
        
        fifo_inputs_140248006750728(0) <= outputs_140248006750784(1);
        outputs_full_140248006750784(1) <= fifo_full_140248006750728(0);
        
        fifo_inputs_140248006750896(1) <= outputs_140248006750840(0);
        outputs_full_140248006750840(0) <= fifo_full_140248006750896(1);
        
        fifo_inputs_140248006750784(0) <= outputs_140248006750840(1);
        outputs_full_140248006750840(1) <= fifo_full_140248006750784(0);
        
        fifo_inputs_140248006750952(1) <= outputs_140248006750896(0);
        outputs_full_140248006750896(0) <= fifo_full_140248006750952(1);
        
        fifo_inputs_140248006750840(0) <= outputs_140248006750896(1);
        outputs_full_140248006750896(1) <= fifo_full_140248006750840(0);
        
        fifo_inputs_140248006751008(1) <= outputs_140248006750952(0);
        outputs_full_140248006750952(0) <= fifo_full_140248006751008(1);
        
        fifo_inputs_140248006750896(0) <= outputs_140248006750952(1);
        outputs_full_140248006750952(1) <= fifo_full_140248006750896(0);
        
        fifo_inputs_140248006751064(1) <= outputs_140248006751008(0);
        outputs_full_140248006751008(0) <= fifo_full_140248006751064(1);
        
        fifo_inputs_140248006750952(0) <= outputs_140248006751008(1);
        outputs_full_140248006751008(1) <= fifo_full_140248006750952(0);
        
        fifo_inputs_140248006751120(1) <= outputs_140248006751064(0);
        outputs_full_140248006751064(0) <= fifo_full_140248006751120(1);
        
        fifo_inputs_140248006751008(0) <= outputs_140248006751064(1);
        outputs_full_140248006751064(1) <= fifo_full_140248006751008(0);
        
        fifo_inputs_140248006751176(1) <= outputs_140248006751120(0);
        outputs_full_140248006751120(0) <= fifo_full_140248006751176(1);
        
        fifo_inputs_140248006751064(0) <= outputs_140248006751120(1);
        outputs_full_140248006751120(1) <= fifo_full_140248006751064(0);
        
        fifo_inputs_140248006751232(1) <= outputs_140248006751176(0);
        outputs_full_140248006751176(0) <= fifo_full_140248006751232(1);
        
        fifo_inputs_140248006751120(0) <= outputs_140248006751176(1);
        outputs_full_140248006751176(1) <= fifo_full_140248006751120(0);
        
        fifo_inputs_140248006751288(1) <= outputs_140248006751232(0);
        outputs_full_140248006751232(0) <= fifo_full_140248006751288(1);
        
        fifo_inputs_140248006751176(0) <= outputs_140248006751232(1);
        outputs_full_140248006751232(1) <= fifo_full_140248006751176(0);
        
        fifo_inputs_140248006751344(1) <= outputs_140248006751288(0);
        outputs_full_140248006751288(0) <= fifo_full_140248006751344(1);
        
        fifo_inputs_140248006751232(0) <= outputs_140248006751288(1);
        outputs_full_140248006751288(1) <= fifo_full_140248006751232(0);
        
        fifo_inputs_140248006751400(1) <= outputs_140248006751344(0);
        outputs_full_140248006751344(0) <= fifo_full_140248006751400(1);
        
        fifo_inputs_140248006751288(0) <= outputs_140248006751344(1);
        outputs_full_140248006751344(1) <= fifo_full_140248006751288(0);
        
        fifo_inputs_140248006751456(1) <= outputs_140248006751400(0);
        outputs_full_140248006751400(0) <= fifo_full_140248006751456(1);
        
        fifo_inputs_140248006751344(0) <= outputs_140248006751400(1);
        outputs_full_140248006751400(1) <= fifo_full_140248006751344(0);
        
        fifo_inputs_140248006751512(1) <= outputs_140248006751456(0);
        outputs_full_140248006751456(0) <= fifo_full_140248006751512(1);
        
        fifo_inputs_140248006751400(0) <= outputs_140248006751456(1);
        outputs_full_140248006751456(1) <= fifo_full_140248006751400(0);
        
        fifo_inputs_140248006751568(1) <= outputs_140248006751512(0);
        outputs_full_140248006751512(0) <= fifo_full_140248006751568(1);
        
        fifo_inputs_140248006751456(0) <= outputs_140248006751512(1);
        outputs_full_140248006751512(1) <= fifo_full_140248006751456(0);
        
        fifo_inputs_140248006751624(1) <= outputs_140248006751568(0);
        outputs_full_140248006751568(0) <= fifo_full_140248006751624(1);
        
        fifo_inputs_140248006751512(0) <= outputs_140248006751568(1);
        outputs_full_140248006751568(1) <= fifo_full_140248006751512(0);
        
        fifo_inputs_140248006751680(1) <= outputs_140248006751624(0);
        outputs_full_140248006751624(0) <= fifo_full_140248006751680(1);
        
        fifo_inputs_140248006751568(0) <= outputs_140248006751624(1);
        outputs_full_140248006751624(1) <= fifo_full_140248006751568(0);
        
        fifo_inputs_140248006751736(1) <= outputs_140248006751680(0);
        outputs_full_140248006751680(0) <= fifo_full_140248006751736(1);
        
        fifo_inputs_140248006751624(0) <= outputs_140248006751680(1);
        outputs_full_140248006751680(1) <= fifo_full_140248006751624(0);
        
        fifo_inputs_140248006751792(1) <= outputs_140248006751736(0);
        outputs_full_140248006751736(0) <= fifo_full_140248006751792(1);
        
        fifo_inputs_140248006751680(0) <= outputs_140248006751736(1);
        outputs_full_140248006751736(1) <= fifo_full_140248006751680(0);
        
        fifo_inputs_140248006751848(1) <= outputs_140248006751792(0);
        outputs_full_140248006751792(0) <= fifo_full_140248006751848(1);
        
        fifo_inputs_140248006751736(0) <= outputs_140248006751792(1);
        outputs_full_140248006751792(1) <= fifo_full_140248006751736(0);
        
        fifo_inputs_140248006751904(1) <= outputs_140248006751848(0);
        outputs_full_140248006751848(0) <= fifo_full_140248006751904(1);
        
        fifo_inputs_140248006751792(0) <= outputs_140248006751848(1);
        outputs_full_140248006751848(1) <= fifo_full_140248006751792(0);
        
        fifo_inputs_140248006751960(1) <= outputs_140248006751904(0);
        outputs_full_140248006751904(0) <= fifo_full_140248006751960(1);
        
        fifo_inputs_140248006751848(0) <= outputs_140248006751904(1);
        outputs_full_140248006751904(1) <= fifo_full_140248006751848(0);
        
        fifo_inputs_140248006752016(1) <= outputs_140248006751960(0);
        outputs_full_140248006751960(0) <= fifo_full_140248006752016(1);
        
        fifo_inputs_140248006751904(0) <= outputs_140248006751960(1);
        outputs_full_140248006751960(1) <= fifo_full_140248006751904(0);
        
        fifo_inputs_140248006752072(1) <= outputs_140248006752016(0);
        outputs_full_140248006752016(0) <= fifo_full_140248006752072(1);
        
        fifo_inputs_140248006751960(0) <= outputs_140248006752016(1);
        outputs_full_140248006752016(1) <= fifo_full_140248006751960(0);
        
        fifo_inputs_140248006752128(1) <= outputs_140248006752072(0);
        outputs_full_140248006752072(0) <= fifo_full_140248006752128(1);
        
        fifo_inputs_140248006752016(0) <= outputs_140248006752072(1);
        outputs_full_140248006752072(1) <= fifo_full_140248006752016(0);
        
        fifo_inputs_140248006752184(1) <= outputs_140248006752128(0);
        outputs_full_140248006752128(0) <= fifo_full_140248006752184(1);
        
        fifo_inputs_140248006752072(0) <= outputs_140248006752128(1);
        outputs_full_140248006752128(1) <= fifo_full_140248006752072(0);
        
        fifo_inputs_140248006752240(1) <= outputs_140248006752184(0);
        outputs_full_140248006752184(0) <= fifo_full_140248006752240(1);
        
        fifo_inputs_140248006752128(0) <= outputs_140248006752184(1);
        outputs_full_140248006752184(1) <= fifo_full_140248006752128(0);
        
        fifo_inputs_140248006752296(1) <= outputs_140248006752240(0);
        outputs_full_140248006752240(0) <= fifo_full_140248006752296(1);
        
        fifo_inputs_140248006752184(0) <= outputs_140248006752240(1);
        outputs_full_140248006752240(1) <= fifo_full_140248006752184(0);
        
        fifo_inputs_140248006752352(1) <= outputs_140248006752296(0);
        outputs_full_140248006752296(0) <= fifo_full_140248006752352(1);
        
        fifo_inputs_140248006752240(0) <= outputs_140248006752296(1);
        outputs_full_140248006752296(1) <= fifo_full_140248006752240(0);
        
        fifo_inputs_140248006752408(1) <= outputs_140248006752352(0);
        outputs_full_140248006752352(0) <= fifo_full_140248006752408(1);
        
        fifo_inputs_140248006752296(0) <= outputs_140248006752352(1);
        outputs_full_140248006752352(1) <= fifo_full_140248006752296(0);
        
        fifo_inputs_140248006752352(0) <= outputs_140248006752408(1);
        outputs_full_140248006752408(1) <= fifo_full_140248006752352(0);
        

    
        core_inst_140248006679688: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006679688,
            fifo_full => fifo_full_140248006679688,
            outputs => outputs_140248006679688,
            outputs_full => outputs_full_140248006679688
        );
        
        core_inst_140248006679632: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006679632,
            fifo_full => fifo_full_140248006679632,
            outputs => outputs_140248006679632,
            outputs_full => outputs_full_140248006679632
        );
        
        core_inst_140248006679856: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006679856,
            fifo_full => fifo_full_140248006679856,
            outputs => outputs_140248006679856,
            outputs_full => outputs_full_140248006679856
        );
        
        core_inst_140248006679912: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006679912,
            fifo_full => fifo_full_140248006679912,
            outputs => outputs_140248006679912,
            outputs_full => outputs_full_140248006679912
        );
        
        core_inst_140248006679968: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006679968,
            fifo_full => fifo_full_140248006679968,
            outputs => outputs_140248006679968,
            outputs_full => outputs_full_140248006679968
        );
        
        core_inst_140248006679800: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006679800,
            fifo_full => fifo_full_140248006679800,
            outputs => outputs_140248006679800,
            outputs_full => outputs_full_140248006679800
        );
        
        core_inst_140248006680024: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006680024,
            fifo_full => fifo_full_140248006680024,
            outputs => outputs_140248006680024,
            outputs_full => outputs_full_140248006680024
        );
        
        core_inst_140248006680080: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006680080,
            fifo_full => fifo_full_140248006680080,
            outputs => outputs_140248006680080,
            outputs_full => outputs_full_140248006680080
        );
        
        core_inst_140248006680136: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006680136,
            fifo_full => fifo_full_140248006680136,
            outputs => outputs_140248006680136,
            outputs_full => outputs_full_140248006680136
        );
        
        core_inst_140248006680192: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006680192,
            fifo_full => fifo_full_140248006680192,
            outputs => outputs_140248006680192,
            outputs_full => outputs_full_140248006680192
        );
        
        core_inst_140248006679744: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006679744,
            fifo_full => fifo_full_140248006679744,
            outputs => outputs_140248006679744,
            outputs_full => outputs_full_140248006679744
        );
        
        core_inst_140248006680248: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006680248,
            fifo_full => fifo_full_140248006680248,
            outputs => outputs_140248006680248,
            outputs_full => outputs_full_140248006680248
        );
        
        core_inst_140248006680304: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006680304,
            fifo_full => fifo_full_140248006680304,
            outputs => outputs_140248006680304,
            outputs_full => outputs_full_140248006680304
        );
        
        core_inst_140248006680360: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006680360,
            fifo_full => fifo_full_140248006680360,
            outputs => outputs_140248006680360,
            outputs_full => outputs_full_140248006680360
        );
        
        core_inst_140248006680416: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006680416,
            fifo_full => fifo_full_140248006680416,
            outputs => outputs_140248006680416,
            outputs_full => outputs_full_140248006680416
        );
        
        core_inst_140248006680472: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006680472,
            fifo_full => fifo_full_140248006680472,
            outputs => outputs_140248006680472,
            outputs_full => outputs_full_140248006680472
        );
        
        core_inst_140248006680528: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006680528,
            fifo_full => fifo_full_140248006680528,
            outputs => outputs_140248006680528,
            outputs_full => outputs_full_140248006680528
        );
        
        core_inst_140248006729800: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006729800,
            fifo_full => fifo_full_140248006729800,
            outputs => outputs_140248006729800,
            outputs_full => outputs_full_140248006729800
        );
        
        core_inst_140248006729856: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006729856,
            fifo_full => fifo_full_140248006729856,
            outputs => outputs_140248006729856,
            outputs_full => outputs_full_140248006729856
        );
        
        core_inst_140248006729912: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006729912,
            fifo_full => fifo_full_140248006729912,
            outputs => outputs_140248006729912,
            outputs_full => outputs_full_140248006729912
        );
        
        core_inst_140248006729968: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006729968,
            fifo_full => fifo_full_140248006729968,
            outputs => outputs_140248006729968,
            outputs_full => outputs_full_140248006729968
        );
        
        core_inst_140248006730024: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006730024,
            fifo_full => fifo_full_140248006730024,
            outputs => outputs_140248006730024,
            outputs_full => outputs_full_140248006730024
        );
        
        core_inst_140248006730080: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006730080,
            fifo_full => fifo_full_140248006730080,
            outputs => outputs_140248006730080,
            outputs_full => outputs_full_140248006730080
        );
        
        core_inst_140248006730136: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006730136,
            fifo_full => fifo_full_140248006730136,
            outputs => outputs_140248006730136,
            outputs_full => outputs_full_140248006730136
        );
        
        core_inst_140248006730192: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006730192,
            fifo_full => fifo_full_140248006730192,
            outputs => outputs_140248006730192,
            outputs_full => outputs_full_140248006730192
        );
        
        core_inst_140248006730248: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006730248,
            fifo_full => fifo_full_140248006730248,
            outputs => outputs_140248006730248,
            outputs_full => outputs_full_140248006730248
        );
        
        core_inst_140248006730304: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006730304,
            fifo_full => fifo_full_140248006730304,
            outputs => outputs_140248006730304,
            outputs_full => outputs_full_140248006730304
        );
        
        core_inst_140248006730360: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006730360,
            fifo_full => fifo_full_140248006730360,
            outputs => outputs_140248006730360,
            outputs_full => outputs_full_140248006730360
        );
        
        core_inst_140248006730416: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006730416,
            fifo_full => fifo_full_140248006730416,
            outputs => outputs_140248006730416,
            outputs_full => outputs_full_140248006730416
        );
        
        core_inst_140248006730472: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006730472,
            fifo_full => fifo_full_140248006730472,
            outputs => outputs_140248006730472,
            outputs_full => outputs_full_140248006730472
        );
        
        core_inst_140248006730528: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006730528,
            fifo_full => fifo_full_140248006730528,
            outputs => outputs_140248006730528,
            outputs_full => outputs_full_140248006730528
        );
        
        core_inst_140248006730584: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006730584,
            fifo_full => fifo_full_140248006730584,
            outputs => outputs_140248006730584,
            outputs_full => outputs_full_140248006730584
        );
        
        core_inst_140248006730640: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006730640,
            fifo_full => fifo_full_140248006730640,
            outputs => outputs_140248006730640,
            outputs_full => outputs_full_140248006730640
        );
        
        core_inst_140248006730696: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006730696,
            fifo_full => fifo_full_140248006730696,
            outputs => outputs_140248006730696,
            outputs_full => outputs_full_140248006730696
        );
        
        core_inst_140248006730752: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006730752,
            fifo_full => fifo_full_140248006730752,
            outputs => outputs_140248006730752,
            outputs_full => outputs_full_140248006730752
        );
        
        core_inst_140248006730808: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006730808,
            fifo_full => fifo_full_140248006730808,
            outputs => outputs_140248006730808,
            outputs_full => outputs_full_140248006730808
        );
        
        core_inst_140248006730864: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006730864,
            fifo_full => fifo_full_140248006730864,
            outputs => outputs_140248006730864,
            outputs_full => outputs_full_140248006730864
        );
        
        core_inst_140248006730920: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006730920,
            fifo_full => fifo_full_140248006730920,
            outputs => outputs_140248006730920,
            outputs_full => outputs_full_140248006730920
        );
        
        core_inst_140248006730976: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006730976,
            fifo_full => fifo_full_140248006730976,
            outputs => outputs_140248006730976,
            outputs_full => outputs_full_140248006730976
        );
        
        core_inst_140248006731032: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006731032,
            fifo_full => fifo_full_140248006731032,
            outputs => outputs_140248006731032,
            outputs_full => outputs_full_140248006731032
        );
        
        core_inst_140248006731088: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006731088,
            fifo_full => fifo_full_140248006731088,
            outputs => outputs_140248006731088,
            outputs_full => outputs_full_140248006731088
        );
        
        core_inst_140248006731144: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006731144,
            fifo_full => fifo_full_140248006731144,
            outputs => outputs_140248006731144,
            outputs_full => outputs_full_140248006731144
        );
        
        core_inst_140248006731200: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006731200,
            fifo_full => fifo_full_140248006731200,
            outputs => outputs_140248006731200,
            outputs_full => outputs_full_140248006731200
        );
        
        core_inst_140248006731256: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006731256,
            fifo_full => fifo_full_140248006731256,
            outputs => outputs_140248006731256,
            outputs_full => outputs_full_140248006731256
        );
        
        core_inst_140248006731312: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006731312,
            fifo_full => fifo_full_140248006731312,
            outputs => outputs_140248006731312,
            outputs_full => outputs_full_140248006731312
        );
        
        core_inst_140248006731368: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006731368,
            fifo_full => fifo_full_140248006731368,
            outputs => outputs_140248006731368,
            outputs_full => outputs_full_140248006731368
        );
        
        core_inst_140248006731424: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006731424,
            fifo_full => fifo_full_140248006731424,
            outputs => outputs_140248006731424,
            outputs_full => outputs_full_140248006731424
        );
        
        core_inst_140248006731480: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006731480,
            fifo_full => fifo_full_140248006731480,
            outputs => outputs_140248006731480,
            outputs_full => outputs_full_140248006731480
        );
        
        core_inst_140248006731536: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006731536,
            fifo_full => fifo_full_140248006731536,
            outputs => outputs_140248006731536,
            outputs_full => outputs_full_140248006731536
        );
        
        core_inst_140248006731592: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006731592,
            fifo_full => fifo_full_140248006731592,
            outputs => outputs_140248006731592,
            outputs_full => outputs_full_140248006731592
        );
        
        core_inst_140248006731648: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006731648,
            fifo_full => fifo_full_140248006731648,
            outputs => outputs_140248006731648,
            outputs_full => outputs_full_140248006731648
        );
        
        core_inst_140248006731704: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006731704,
            fifo_full => fifo_full_140248006731704,
            outputs => outputs_140248006731704,
            outputs_full => outputs_full_140248006731704
        );
        
        core_inst_140248006731760: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006731760,
            fifo_full => fifo_full_140248006731760,
            outputs => outputs_140248006731760,
            outputs_full => outputs_full_140248006731760
        );
        
        core_inst_140248006731816: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006731816,
            fifo_full => fifo_full_140248006731816,
            outputs => outputs_140248006731816,
            outputs_full => outputs_full_140248006731816
        );
        
        core_inst_140248006731872: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006731872,
            fifo_full => fifo_full_140248006731872,
            outputs => outputs_140248006731872,
            outputs_full => outputs_full_140248006731872
        );
        
        core_inst_140248006731928: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006731928,
            fifo_full => fifo_full_140248006731928,
            outputs => outputs_140248006731928,
            outputs_full => outputs_full_140248006731928
        );
        
        core_inst_140248006731984: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006731984,
            fifo_full => fifo_full_140248006731984,
            outputs => outputs_140248006731984,
            outputs_full => outputs_full_140248006731984
        );
        
        core_inst_140248006732040: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006732040,
            fifo_full => fifo_full_140248006732040,
            outputs => outputs_140248006732040,
            outputs_full => outputs_full_140248006732040
        );
        
        core_inst_140248006732096: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006732096,
            fifo_full => fifo_full_140248006732096,
            outputs => outputs_140248006732096,
            outputs_full => outputs_full_140248006732096
        );
        
        core_inst_140248006732152: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006732152,
            fifo_full => fifo_full_140248006732152,
            outputs => outputs_140248006732152,
            outputs_full => outputs_full_140248006732152
        );
        
        core_inst_140248006732208: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006732208,
            fifo_full => fifo_full_140248006732208,
            outputs => outputs_140248006732208,
            outputs_full => outputs_full_140248006732208
        );
        
        core_inst_140248006732264: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006732264,
            fifo_full => fifo_full_140248006732264,
            outputs => outputs_140248006732264,
            outputs_full => outputs_full_140248006732264
        );
        
        core_inst_140248006732320: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006732320,
            fifo_full => fifo_full_140248006732320,
            outputs => outputs_140248006732320,
            outputs_full => outputs_full_140248006732320
        );
        
        core_inst_140248006732376: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006732376,
            fifo_full => fifo_full_140248006732376,
            outputs => outputs_140248006732376,
            outputs_full => outputs_full_140248006732376
        );
        
        core_inst_140248006732432: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006732432,
            fifo_full => fifo_full_140248006732432,
            outputs => outputs_140248006732432,
            outputs_full => outputs_full_140248006732432
        );
        
        core_inst_140248006732488: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006732488,
            fifo_full => fifo_full_140248006732488,
            outputs => outputs_140248006732488,
            outputs_full => outputs_full_140248006732488
        );
        
        core_inst_140248006732544: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006732544,
            fifo_full => fifo_full_140248006732544,
            outputs => outputs_140248006732544,
            outputs_full => outputs_full_140248006732544
        );
        
        core_inst_140248006732600: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006732600,
            fifo_full => fifo_full_140248006732600,
            outputs => outputs_140248006732600,
            outputs_full => outputs_full_140248006732600
        );
        
        core_inst_140248006732656: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006732656,
            fifo_full => fifo_full_140248006732656,
            outputs => outputs_140248006732656,
            outputs_full => outputs_full_140248006732656
        );
        
        core_inst_140248006732712: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006732712,
            fifo_full => fifo_full_140248006732712,
            outputs => outputs_140248006732712,
            outputs_full => outputs_full_140248006732712
        );
        
        core_inst_140248006732768: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006732768,
            fifo_full => fifo_full_140248006732768,
            outputs => outputs_140248006732768,
            outputs_full => outputs_full_140248006732768
        );
        
        core_inst_140248006732824: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006732824,
            fifo_full => fifo_full_140248006732824,
            outputs => outputs_140248006732824,
            outputs_full => outputs_full_140248006732824
        );
        
        core_inst_140248006732880: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006732880,
            fifo_full => fifo_full_140248006732880,
            outputs => outputs_140248006732880,
            outputs_full => outputs_full_140248006732880
        );
        
        core_inst_140248006732936: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006732936,
            fifo_full => fifo_full_140248006732936,
            outputs => outputs_140248006732936,
            outputs_full => outputs_full_140248006732936
        );
        
        core_inst_140248006732992: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006732992,
            fifo_full => fifo_full_140248006732992,
            outputs => outputs_140248006732992,
            outputs_full => outputs_full_140248006732992
        );
        
        core_inst_140248006733048: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006733048,
            fifo_full => fifo_full_140248006733048,
            outputs => outputs_140248006733048,
            outputs_full => outputs_full_140248006733048
        );
        
        core_inst_140248006733104: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006733104,
            fifo_full => fifo_full_140248006733104,
            outputs => outputs_140248006733104,
            outputs_full => outputs_full_140248006733104
        );
        
        core_inst_140248006733160: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006733160,
            fifo_full => fifo_full_140248006733160,
            outputs => outputs_140248006733160,
            outputs_full => outputs_full_140248006733160
        );
        
        core_inst_140248006733216: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006733216,
            fifo_full => fifo_full_140248006733216,
            outputs => outputs_140248006733216,
            outputs_full => outputs_full_140248006733216
        );
        
        core_inst_140248006733272: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006733272,
            fifo_full => fifo_full_140248006733272,
            outputs => outputs_140248006733272,
            outputs_full => outputs_full_140248006733272
        );
        
        core_inst_140248006733328: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006733328,
            fifo_full => fifo_full_140248006733328,
            outputs => outputs_140248006733328,
            outputs_full => outputs_full_140248006733328
        );
        
        core_inst_140248006733384: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006733384,
            fifo_full => fifo_full_140248006733384,
            outputs => outputs_140248006733384,
            outputs_full => outputs_full_140248006733384
        );
        
        core_inst_140248006733440: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006733440,
            fifo_full => fifo_full_140248006733440,
            outputs => outputs_140248006733440,
            outputs_full => outputs_full_140248006733440
        );
        
        core_inst_140248006733496: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006733496,
            fifo_full => fifo_full_140248006733496,
            outputs => outputs_140248006733496,
            outputs_full => outputs_full_140248006733496
        );
        
        core_inst_140248006733552: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006733552,
            fifo_full => fifo_full_140248006733552,
            outputs => outputs_140248006733552,
            outputs_full => outputs_full_140248006733552
        );
        
        core_inst_140248006733608: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006733608,
            fifo_full => fifo_full_140248006733608,
            outputs => outputs_140248006733608,
            outputs_full => outputs_full_140248006733608
        );
        
        core_inst_140248006733664: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006733664,
            fifo_full => fifo_full_140248006733664,
            outputs => outputs_140248006733664,
            outputs_full => outputs_full_140248006733664
        );
        
        core_inst_140248006733720: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006733720,
            fifo_full => fifo_full_140248006733720,
            outputs => outputs_140248006733720,
            outputs_full => outputs_full_140248006733720
        );
        
        core_inst_140248006733776: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006733776,
            fifo_full => fifo_full_140248006733776,
            outputs => outputs_140248006733776,
            outputs_full => outputs_full_140248006733776
        );
        
        core_inst_140248006750280: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006750280,
            fifo_full => fifo_full_140248006750280,
            outputs => outputs_140248006750280,
            outputs_full => outputs_full_140248006750280
        );
        
        core_inst_140248006750336: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006750336,
            fifo_full => fifo_full_140248006750336,
            outputs => outputs_140248006750336,
            outputs_full => outputs_full_140248006750336
        );
        
        core_inst_140248006750392: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006750392,
            fifo_full => fifo_full_140248006750392,
            outputs => outputs_140248006750392,
            outputs_full => outputs_full_140248006750392
        );
        
        core_inst_140248006750448: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006750448,
            fifo_full => fifo_full_140248006750448,
            outputs => outputs_140248006750448,
            outputs_full => outputs_full_140248006750448
        );
        
        core_inst_140248006750504: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006750504,
            fifo_full => fifo_full_140248006750504,
            outputs => outputs_140248006750504,
            outputs_full => outputs_full_140248006750504
        );
        
        core_inst_140248006750560: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006750560,
            fifo_full => fifo_full_140248006750560,
            outputs => outputs_140248006750560,
            outputs_full => outputs_full_140248006750560
        );
        
        core_inst_140248006750616: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006750616,
            fifo_full => fifo_full_140248006750616,
            outputs => outputs_140248006750616,
            outputs_full => outputs_full_140248006750616
        );
        
        core_inst_140248006750672: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006750672,
            fifo_full => fifo_full_140248006750672,
            outputs => outputs_140248006750672,
            outputs_full => outputs_full_140248006750672
        );
        
        core_inst_140248006750728: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006750728,
            fifo_full => fifo_full_140248006750728,
            outputs => outputs_140248006750728,
            outputs_full => outputs_full_140248006750728
        );
        
        core_inst_140248006750784: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006750784,
            fifo_full => fifo_full_140248006750784,
            outputs => outputs_140248006750784,
            outputs_full => outputs_full_140248006750784
        );
        
        core_inst_140248006750840: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006750840,
            fifo_full => fifo_full_140248006750840,
            outputs => outputs_140248006750840,
            outputs_full => outputs_full_140248006750840
        );
        
        core_inst_140248006750896: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006750896,
            fifo_full => fifo_full_140248006750896,
            outputs => outputs_140248006750896,
            outputs_full => outputs_full_140248006750896
        );
        
        core_inst_140248006750952: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006750952,
            fifo_full => fifo_full_140248006750952,
            outputs => outputs_140248006750952,
            outputs_full => outputs_full_140248006750952
        );
        
        core_inst_140248006751008: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006751008,
            fifo_full => fifo_full_140248006751008,
            outputs => outputs_140248006751008,
            outputs_full => outputs_full_140248006751008
        );
        
        core_inst_140248006751064: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006751064,
            fifo_full => fifo_full_140248006751064,
            outputs => outputs_140248006751064,
            outputs_full => outputs_full_140248006751064
        );
        
        core_inst_140248006751120: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006751120,
            fifo_full => fifo_full_140248006751120,
            outputs => outputs_140248006751120,
            outputs_full => outputs_full_140248006751120
        );
        
        core_inst_140248006751176: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006751176,
            fifo_full => fifo_full_140248006751176,
            outputs => outputs_140248006751176,
            outputs_full => outputs_full_140248006751176
        );
        
        core_inst_140248006751232: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006751232,
            fifo_full => fifo_full_140248006751232,
            outputs => outputs_140248006751232,
            outputs_full => outputs_full_140248006751232
        );
        
        core_inst_140248006751288: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006751288,
            fifo_full => fifo_full_140248006751288,
            outputs => outputs_140248006751288,
            outputs_full => outputs_full_140248006751288
        );
        
        core_inst_140248006751344: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006751344,
            fifo_full => fifo_full_140248006751344,
            outputs => outputs_140248006751344,
            outputs_full => outputs_full_140248006751344
        );
        
        core_inst_140248006751400: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006751400,
            fifo_full => fifo_full_140248006751400,
            outputs => outputs_140248006751400,
            outputs_full => outputs_full_140248006751400
        );
        
        core_inst_140248006751456: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006751456,
            fifo_full => fifo_full_140248006751456,
            outputs => outputs_140248006751456,
            outputs_full => outputs_full_140248006751456
        );
        
        core_inst_140248006751512: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006751512,
            fifo_full => fifo_full_140248006751512,
            outputs => outputs_140248006751512,
            outputs_full => outputs_full_140248006751512
        );
        
        core_inst_140248006751568: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006751568,
            fifo_full => fifo_full_140248006751568,
            outputs => outputs_140248006751568,
            outputs_full => outputs_full_140248006751568
        );
        
        core_inst_140248006751624: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006751624,
            fifo_full => fifo_full_140248006751624,
            outputs => outputs_140248006751624,
            outputs_full => outputs_full_140248006751624
        );
        
        core_inst_140248006751680: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006751680,
            fifo_full => fifo_full_140248006751680,
            outputs => outputs_140248006751680,
            outputs_full => outputs_full_140248006751680
        );
        
        core_inst_140248006751736: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006751736,
            fifo_full => fifo_full_140248006751736,
            outputs => outputs_140248006751736,
            outputs_full => outputs_full_140248006751736
        );
        
        core_inst_140248006751792: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006751792,
            fifo_full => fifo_full_140248006751792,
            outputs => outputs_140248006751792,
            outputs_full => outputs_full_140248006751792
        );
        
        core_inst_140248006751848: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006751848,
            fifo_full => fifo_full_140248006751848,
            outputs => outputs_140248006751848,
            outputs_full => outputs_full_140248006751848
        );
        
        core_inst_140248006751904: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006751904,
            fifo_full => fifo_full_140248006751904,
            outputs => outputs_140248006751904,
            outputs_full => outputs_full_140248006751904
        );
        
        core_inst_140248006751960: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006751960,
            fifo_full => fifo_full_140248006751960,
            outputs => outputs_140248006751960,
            outputs_full => outputs_full_140248006751960
        );
        
        core_inst_140248006752016: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006752016,
            fifo_full => fifo_full_140248006752016,
            outputs => outputs_140248006752016,
            outputs_full => outputs_full_140248006752016
        );
        
        core_inst_140248006752072: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006752072,
            fifo_full => fifo_full_140248006752072,
            outputs => outputs_140248006752072,
            outputs_full => outputs_full_140248006752072
        );
        
        core_inst_140248006752128: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006752128,
            fifo_full => fifo_full_140248006752128,
            outputs => outputs_140248006752128,
            outputs_full => outputs_full_140248006752128
        );
        
        core_inst_140248006752184: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006752184,
            fifo_full => fifo_full_140248006752184,
            outputs => outputs_140248006752184,
            outputs_full => outputs_full_140248006752184
        );
        
        core_inst_140248006752240: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006752240,
            fifo_full => fifo_full_140248006752240,
            outputs => outputs_140248006752240,
            outputs_full => outputs_full_140248006752240
        );
        
        core_inst_140248006752296: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006752296,
            fifo_full => fifo_full_140248006752296,
            outputs => outputs_140248006752296,
            outputs_full => outputs_full_140248006752296
        );
        
        core_inst_140248006752352: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006752352,
            fifo_full => fifo_full_140248006752352,
            outputs => outputs_140248006752352,
            outputs_full => outputs_full_140248006752352
        );
        
        core_inst_140248006752408: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_140248006752408,
            fifo_full => fifo_full_140248006752408,
            outputs => outputs_140248006752408,
            outputs_full => outputs_full_140248006752408
        );
        

end behav;

