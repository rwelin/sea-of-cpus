library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity Core is
    port (
        clk: std_logic
    );
end Core;

architecture behav of Core is

begin


end behav;
