
library ieee;
use ieee.std_logic_1164.all;
use work.core_config.all;
use work.all;

entity Grid8x8 is
    port (
        clk: in std_logic;
        clk_en: in std_logic;
        reset: in std_logic;
        addr: in ram_addr;
        data: in word;
        we: in std_logic;
        fifo_inputs: in core_fifo_inputs_t;
        fifo_full: out std_logic_vector(0 to NUM_CORE_FIFOS-1);
        outputs: out core_fifo_inputs_t;
        outputs_full: in std_logic_vector(0 to NUM_CORE_FIFOS-1)
    );
end Grid8x8;

architecture behav of Grid8x8 is

    
        signal fifo_inputs_139867185248632: core_fifo_inputs_t;
        signal fifo_full_139867185248632: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185248632: core_fifo_inputs_t;
        signal outputs_full_139867185248632: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185248856: core_fifo_inputs_t;
        signal fifo_full_139867185248856: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185248856: core_fifo_inputs_t;
        signal outputs_full_139867185248856: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185248912: core_fifo_inputs_t;
        signal fifo_full_139867185248912: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185248912: core_fifo_inputs_t;
        signal outputs_full_139867185248912: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185248968: core_fifo_inputs_t;
        signal fifo_full_139867185248968: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185248968: core_fifo_inputs_t;
        signal outputs_full_139867185248968: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185248800: core_fifo_inputs_t;
        signal fifo_full_139867185248800: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185248800: core_fifo_inputs_t;
        signal outputs_full_139867185248800: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185249024: core_fifo_inputs_t;
        signal fifo_full_139867185249024: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185249024: core_fifo_inputs_t;
        signal outputs_full_139867185249024: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185249080: core_fifo_inputs_t;
        signal fifo_full_139867185249080: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185249080: core_fifo_inputs_t;
        signal outputs_full_139867185249080: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185249136: core_fifo_inputs_t;
        signal fifo_full_139867185249136: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185249136: core_fifo_inputs_t;
        signal outputs_full_139867185249136: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185249192: core_fifo_inputs_t;
        signal fifo_full_139867185249192: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185249192: core_fifo_inputs_t;
        signal outputs_full_139867185249192: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185248744: core_fifo_inputs_t;
        signal fifo_full_139867185248744: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185248744: core_fifo_inputs_t;
        signal outputs_full_139867185248744: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185249248: core_fifo_inputs_t;
        signal fifo_full_139867185249248: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185249248: core_fifo_inputs_t;
        signal outputs_full_139867185249248: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185249304: core_fifo_inputs_t;
        signal fifo_full_139867185249304: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185249304: core_fifo_inputs_t;
        signal outputs_full_139867185249304: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185249360: core_fifo_inputs_t;
        signal fifo_full_139867185249360: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185249360: core_fifo_inputs_t;
        signal outputs_full_139867185249360: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185249416: core_fifo_inputs_t;
        signal fifo_full_139867185249416: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185249416: core_fifo_inputs_t;
        signal outputs_full_139867185249416: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185249472: core_fifo_inputs_t;
        signal fifo_full_139867185249472: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185249472: core_fifo_inputs_t;
        signal outputs_full_139867185249472: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185249528: core_fifo_inputs_t;
        signal fifo_full_139867185249528: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185249528: core_fifo_inputs_t;
        signal outputs_full_139867185249528: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185249584: core_fifo_inputs_t;
        signal fifo_full_139867185249584: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185249584: core_fifo_inputs_t;
        signal outputs_full_139867185249584: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185249640: core_fifo_inputs_t;
        signal fifo_full_139867185249640: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185249640: core_fifo_inputs_t;
        signal outputs_full_139867185249640: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185249696: core_fifo_inputs_t;
        signal fifo_full_139867185249696: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185249696: core_fifo_inputs_t;
        signal outputs_full_139867185249696: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185249752: core_fifo_inputs_t;
        signal fifo_full_139867185249752: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185249752: core_fifo_inputs_t;
        signal outputs_full_139867185249752: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185249808: core_fifo_inputs_t;
        signal fifo_full_139867185249808: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185249808: core_fifo_inputs_t;
        signal outputs_full_139867185249808: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185249864: core_fifo_inputs_t;
        signal fifo_full_139867185249864: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185249864: core_fifo_inputs_t;
        signal outputs_full_139867185249864: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185249920: core_fifo_inputs_t;
        signal fifo_full_139867185249920: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185249920: core_fifo_inputs_t;
        signal outputs_full_139867185249920: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185249976: core_fifo_inputs_t;
        signal fifo_full_139867185249976: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185249976: core_fifo_inputs_t;
        signal outputs_full_139867185249976: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185250032: core_fifo_inputs_t;
        signal fifo_full_139867185250032: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185250032: core_fifo_inputs_t;
        signal outputs_full_139867185250032: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185250088: core_fifo_inputs_t;
        signal fifo_full_139867185250088: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185250088: core_fifo_inputs_t;
        signal outputs_full_139867185250088: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185250144: core_fifo_inputs_t;
        signal fifo_full_139867185250144: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185250144: core_fifo_inputs_t;
        signal outputs_full_139867185250144: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185250200: core_fifo_inputs_t;
        signal fifo_full_139867185250200: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185250200: core_fifo_inputs_t;
        signal outputs_full_139867185250200: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185250256: core_fifo_inputs_t;
        signal fifo_full_139867185250256: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185250256: core_fifo_inputs_t;
        signal outputs_full_139867185250256: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185291336: core_fifo_inputs_t;
        signal fifo_full_139867185291336: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185291336: core_fifo_inputs_t;
        signal outputs_full_139867185291336: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185291392: core_fifo_inputs_t;
        signal fifo_full_139867185291392: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185291392: core_fifo_inputs_t;
        signal outputs_full_139867185291392: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185291448: core_fifo_inputs_t;
        signal fifo_full_139867185291448: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185291448: core_fifo_inputs_t;
        signal outputs_full_139867185291448: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185291504: core_fifo_inputs_t;
        signal fifo_full_139867185291504: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185291504: core_fifo_inputs_t;
        signal outputs_full_139867185291504: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185291560: core_fifo_inputs_t;
        signal fifo_full_139867185291560: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185291560: core_fifo_inputs_t;
        signal outputs_full_139867185291560: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185291616: core_fifo_inputs_t;
        signal fifo_full_139867185291616: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185291616: core_fifo_inputs_t;
        signal outputs_full_139867185291616: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185291672: core_fifo_inputs_t;
        signal fifo_full_139867185291672: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185291672: core_fifo_inputs_t;
        signal outputs_full_139867185291672: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185291728: core_fifo_inputs_t;
        signal fifo_full_139867185291728: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185291728: core_fifo_inputs_t;
        signal outputs_full_139867185291728: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185291784: core_fifo_inputs_t;
        signal fifo_full_139867185291784: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185291784: core_fifo_inputs_t;
        signal outputs_full_139867185291784: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185291840: core_fifo_inputs_t;
        signal fifo_full_139867185291840: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185291840: core_fifo_inputs_t;
        signal outputs_full_139867185291840: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185291896: core_fifo_inputs_t;
        signal fifo_full_139867185291896: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185291896: core_fifo_inputs_t;
        signal outputs_full_139867185291896: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185291952: core_fifo_inputs_t;
        signal fifo_full_139867185291952: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185291952: core_fifo_inputs_t;
        signal outputs_full_139867185291952: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185292008: core_fifo_inputs_t;
        signal fifo_full_139867185292008: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185292008: core_fifo_inputs_t;
        signal outputs_full_139867185292008: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185292064: core_fifo_inputs_t;
        signal fifo_full_139867185292064: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185292064: core_fifo_inputs_t;
        signal outputs_full_139867185292064: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185292120: core_fifo_inputs_t;
        signal fifo_full_139867185292120: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185292120: core_fifo_inputs_t;
        signal outputs_full_139867185292120: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185292176: core_fifo_inputs_t;
        signal fifo_full_139867185292176: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185292176: core_fifo_inputs_t;
        signal outputs_full_139867185292176: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185292232: core_fifo_inputs_t;
        signal fifo_full_139867185292232: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185292232: core_fifo_inputs_t;
        signal outputs_full_139867185292232: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185292288: core_fifo_inputs_t;
        signal fifo_full_139867185292288: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185292288: core_fifo_inputs_t;
        signal outputs_full_139867185292288: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185292344: core_fifo_inputs_t;
        signal fifo_full_139867185292344: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185292344: core_fifo_inputs_t;
        signal outputs_full_139867185292344: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185292400: core_fifo_inputs_t;
        signal fifo_full_139867185292400: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185292400: core_fifo_inputs_t;
        signal outputs_full_139867185292400: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185292456: core_fifo_inputs_t;
        signal fifo_full_139867185292456: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185292456: core_fifo_inputs_t;
        signal outputs_full_139867185292456: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185292512: core_fifo_inputs_t;
        signal fifo_full_139867185292512: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185292512: core_fifo_inputs_t;
        signal outputs_full_139867185292512: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185292568: core_fifo_inputs_t;
        signal fifo_full_139867185292568: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185292568: core_fifo_inputs_t;
        signal outputs_full_139867185292568: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185292624: core_fifo_inputs_t;
        signal fifo_full_139867185292624: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185292624: core_fifo_inputs_t;
        signal outputs_full_139867185292624: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185292680: core_fifo_inputs_t;
        signal fifo_full_139867185292680: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185292680: core_fifo_inputs_t;
        signal outputs_full_139867185292680: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185292736: core_fifo_inputs_t;
        signal fifo_full_139867185292736: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185292736: core_fifo_inputs_t;
        signal outputs_full_139867185292736: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185292792: core_fifo_inputs_t;
        signal fifo_full_139867185292792: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185292792: core_fifo_inputs_t;
        signal outputs_full_139867185292792: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185292848: core_fifo_inputs_t;
        signal fifo_full_139867185292848: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185292848: core_fifo_inputs_t;
        signal outputs_full_139867185292848: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185292904: core_fifo_inputs_t;
        signal fifo_full_139867185292904: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185292904: core_fifo_inputs_t;
        signal outputs_full_139867185292904: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185292960: core_fifo_inputs_t;
        signal fifo_full_139867185292960: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185292960: core_fifo_inputs_t;
        signal outputs_full_139867185292960: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185293016: core_fifo_inputs_t;
        signal fifo_full_139867185293016: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185293016: core_fifo_inputs_t;
        signal outputs_full_139867185293016: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185293072: core_fifo_inputs_t;
        signal fifo_full_139867185293072: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185293072: core_fifo_inputs_t;
        signal outputs_full_139867185293072: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185293128: core_fifo_inputs_t;
        signal fifo_full_139867185293128: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185293128: core_fifo_inputs_t;
        signal outputs_full_139867185293128: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185293184: core_fifo_inputs_t;
        signal fifo_full_139867185293184: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185293184: core_fifo_inputs_t;
        signal outputs_full_139867185293184: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        
        signal fifo_inputs_139867185293240: core_fifo_inputs_t;
        signal fifo_full_139867185293240: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        signal outputs_139867185293240: core_fifo_inputs_t;
        signal outputs_full_139867185293240: std_logic_vector(0 to NUM_CORE_FIFOS-1);
        

begin

        outputs(1) <= outputs_139867185248632(1);
        outputs(3) <= outputs_139867185248632(3);
        outputs_full_139867185248632(1) <= outputs_full(1);
        outputs_full_139867185248632(3) <= outputs_full(3);

        outputs(0) <= outputs_139867185293240(0);
        outputs(2) <= outputs_139867185293240(2);
        outputs_full_139867185293240(0) <= outputs_full(0); 
        outputs_full_139867185293240(2) <= outputs_full(2);
    
        fifo_inputs_139867185248856(1) <= outputs_139867185248632(0);
        outputs_full_139867185248632(0) <= fifo_full_139867185248856(1);
        
        fifo_inputs_139867185249192(3) <= outputs_139867185248632(2);
        outputs_full_139867185248632(2) <= fifo_full_139867185249192(3);
        
        fifo_inputs_139867185248912(1) <= outputs_139867185248856(0);
        outputs_full_139867185248856(0) <= fifo_full_139867185248912(1);
        
        fifo_inputs_139867185248632(0) <= outputs_139867185248856(1);
        outputs_full_139867185248856(1) <= fifo_full_139867185248632(0);
        
        fifo_inputs_139867185248744(3) <= outputs_139867185248856(2);
        outputs_full_139867185248856(2) <= fifo_full_139867185248744(3);
        
        fifo_inputs_139867185248968(1) <= outputs_139867185248912(0);
        outputs_full_139867185248912(0) <= fifo_full_139867185248968(1);
        
        fifo_inputs_139867185248856(0) <= outputs_139867185248912(1);
        outputs_full_139867185248912(1) <= fifo_full_139867185248856(0);
        
        fifo_inputs_139867185249248(3) <= outputs_139867185248912(2);
        outputs_full_139867185248912(2) <= fifo_full_139867185249248(3);
        
        fifo_inputs_139867185248800(1) <= outputs_139867185248968(0);
        outputs_full_139867185248968(0) <= fifo_full_139867185248800(1);
        
        fifo_inputs_139867185248912(0) <= outputs_139867185248968(1);
        outputs_full_139867185248968(1) <= fifo_full_139867185248912(0);
        
        fifo_inputs_139867185249304(3) <= outputs_139867185248968(2);
        outputs_full_139867185248968(2) <= fifo_full_139867185249304(3);
        
        fifo_inputs_139867185249024(1) <= outputs_139867185248800(0);
        outputs_full_139867185248800(0) <= fifo_full_139867185249024(1);
        
        fifo_inputs_139867185248968(0) <= outputs_139867185248800(1);
        outputs_full_139867185248800(1) <= fifo_full_139867185248968(0);
        
        fifo_inputs_139867185249360(3) <= outputs_139867185248800(2);
        outputs_full_139867185248800(2) <= fifo_full_139867185249360(3);
        
        fifo_inputs_139867185249080(1) <= outputs_139867185249024(0);
        outputs_full_139867185249024(0) <= fifo_full_139867185249080(1);
        
        fifo_inputs_139867185248800(0) <= outputs_139867185249024(1);
        outputs_full_139867185249024(1) <= fifo_full_139867185248800(0);
        
        fifo_inputs_139867185249416(3) <= outputs_139867185249024(2);
        outputs_full_139867185249024(2) <= fifo_full_139867185249416(3);
        
        fifo_inputs_139867185249136(1) <= outputs_139867185249080(0);
        outputs_full_139867185249080(0) <= fifo_full_139867185249136(1);
        
        fifo_inputs_139867185249024(0) <= outputs_139867185249080(1);
        outputs_full_139867185249080(1) <= fifo_full_139867185249024(0);
        
        fifo_inputs_139867185249472(3) <= outputs_139867185249080(2);
        outputs_full_139867185249080(2) <= fifo_full_139867185249472(3);
        
        fifo_inputs_139867185249080(0) <= outputs_139867185249136(1);
        outputs_full_139867185249136(1) <= fifo_full_139867185249080(0);
        
        fifo_inputs_139867185249528(3) <= outputs_139867185249136(2);
        outputs_full_139867185249136(2) <= fifo_full_139867185249528(3);
        
        fifo_inputs_139867185248744(1) <= outputs_139867185249192(0);
        outputs_full_139867185249192(0) <= fifo_full_139867185248744(1);
        
        fifo_inputs_139867185249584(3) <= outputs_139867185249192(2);
        outputs_full_139867185249192(2) <= fifo_full_139867185249584(3);
        
        fifo_inputs_139867185248632(2) <= outputs_139867185249192(3);
        outputs_full_139867185249192(3) <= fifo_full_139867185248632(2);
        
        fifo_inputs_139867185249248(1) <= outputs_139867185248744(0);
        outputs_full_139867185248744(0) <= fifo_full_139867185249248(1);
        
        fifo_inputs_139867185249192(0) <= outputs_139867185248744(1);
        outputs_full_139867185248744(1) <= fifo_full_139867185249192(0);
        
        fifo_inputs_139867185249640(3) <= outputs_139867185248744(2);
        outputs_full_139867185248744(2) <= fifo_full_139867185249640(3);
        
        fifo_inputs_139867185248856(2) <= outputs_139867185248744(3);
        outputs_full_139867185248744(3) <= fifo_full_139867185248856(2);
        
        fifo_inputs_139867185249304(1) <= outputs_139867185249248(0);
        outputs_full_139867185249248(0) <= fifo_full_139867185249304(1);
        
        fifo_inputs_139867185248744(0) <= outputs_139867185249248(1);
        outputs_full_139867185249248(1) <= fifo_full_139867185248744(0);
        
        fifo_inputs_139867185249696(3) <= outputs_139867185249248(2);
        outputs_full_139867185249248(2) <= fifo_full_139867185249696(3);
        
        fifo_inputs_139867185248912(2) <= outputs_139867185249248(3);
        outputs_full_139867185249248(3) <= fifo_full_139867185248912(2);
        
        fifo_inputs_139867185249360(1) <= outputs_139867185249304(0);
        outputs_full_139867185249304(0) <= fifo_full_139867185249360(1);
        
        fifo_inputs_139867185249248(0) <= outputs_139867185249304(1);
        outputs_full_139867185249304(1) <= fifo_full_139867185249248(0);
        
        fifo_inputs_139867185249752(3) <= outputs_139867185249304(2);
        outputs_full_139867185249304(2) <= fifo_full_139867185249752(3);
        
        fifo_inputs_139867185248968(2) <= outputs_139867185249304(3);
        outputs_full_139867185249304(3) <= fifo_full_139867185248968(2);
        
        fifo_inputs_139867185249416(1) <= outputs_139867185249360(0);
        outputs_full_139867185249360(0) <= fifo_full_139867185249416(1);
        
        fifo_inputs_139867185249304(0) <= outputs_139867185249360(1);
        outputs_full_139867185249360(1) <= fifo_full_139867185249304(0);
        
        fifo_inputs_139867185249808(3) <= outputs_139867185249360(2);
        outputs_full_139867185249360(2) <= fifo_full_139867185249808(3);
        
        fifo_inputs_139867185248800(2) <= outputs_139867185249360(3);
        outputs_full_139867185249360(3) <= fifo_full_139867185248800(2);
        
        fifo_inputs_139867185249472(1) <= outputs_139867185249416(0);
        outputs_full_139867185249416(0) <= fifo_full_139867185249472(1);
        
        fifo_inputs_139867185249360(0) <= outputs_139867185249416(1);
        outputs_full_139867185249416(1) <= fifo_full_139867185249360(0);
        
        fifo_inputs_139867185249864(3) <= outputs_139867185249416(2);
        outputs_full_139867185249416(2) <= fifo_full_139867185249864(3);
        
        fifo_inputs_139867185249024(2) <= outputs_139867185249416(3);
        outputs_full_139867185249416(3) <= fifo_full_139867185249024(2);
        
        fifo_inputs_139867185249528(1) <= outputs_139867185249472(0);
        outputs_full_139867185249472(0) <= fifo_full_139867185249528(1);
        
        fifo_inputs_139867185249416(0) <= outputs_139867185249472(1);
        outputs_full_139867185249472(1) <= fifo_full_139867185249416(0);
        
        fifo_inputs_139867185249920(3) <= outputs_139867185249472(2);
        outputs_full_139867185249472(2) <= fifo_full_139867185249920(3);
        
        fifo_inputs_139867185249080(2) <= outputs_139867185249472(3);
        outputs_full_139867185249472(3) <= fifo_full_139867185249080(2);
        
        fifo_inputs_139867185249472(0) <= outputs_139867185249528(1);
        outputs_full_139867185249528(1) <= fifo_full_139867185249472(0);
        
        fifo_inputs_139867185249976(3) <= outputs_139867185249528(2);
        outputs_full_139867185249528(2) <= fifo_full_139867185249976(3);
        
        fifo_inputs_139867185249136(2) <= outputs_139867185249528(3);
        outputs_full_139867185249528(3) <= fifo_full_139867185249136(2);
        
        fifo_inputs_139867185249640(1) <= outputs_139867185249584(0);
        outputs_full_139867185249584(0) <= fifo_full_139867185249640(1);
        
        fifo_inputs_139867185250032(3) <= outputs_139867185249584(2);
        outputs_full_139867185249584(2) <= fifo_full_139867185250032(3);
        
        fifo_inputs_139867185249192(2) <= outputs_139867185249584(3);
        outputs_full_139867185249584(3) <= fifo_full_139867185249192(2);
        
        fifo_inputs_139867185249696(1) <= outputs_139867185249640(0);
        outputs_full_139867185249640(0) <= fifo_full_139867185249696(1);
        
        fifo_inputs_139867185249584(0) <= outputs_139867185249640(1);
        outputs_full_139867185249640(1) <= fifo_full_139867185249584(0);
        
        fifo_inputs_139867185250088(3) <= outputs_139867185249640(2);
        outputs_full_139867185249640(2) <= fifo_full_139867185250088(3);
        
        fifo_inputs_139867185248744(2) <= outputs_139867185249640(3);
        outputs_full_139867185249640(3) <= fifo_full_139867185248744(2);
        
        fifo_inputs_139867185249752(1) <= outputs_139867185249696(0);
        outputs_full_139867185249696(0) <= fifo_full_139867185249752(1);
        
        fifo_inputs_139867185249640(0) <= outputs_139867185249696(1);
        outputs_full_139867185249696(1) <= fifo_full_139867185249640(0);
        
        fifo_inputs_139867185250144(3) <= outputs_139867185249696(2);
        outputs_full_139867185249696(2) <= fifo_full_139867185250144(3);
        
        fifo_inputs_139867185249248(2) <= outputs_139867185249696(3);
        outputs_full_139867185249696(3) <= fifo_full_139867185249248(2);
        
        fifo_inputs_139867185249808(1) <= outputs_139867185249752(0);
        outputs_full_139867185249752(0) <= fifo_full_139867185249808(1);
        
        fifo_inputs_139867185249696(0) <= outputs_139867185249752(1);
        outputs_full_139867185249752(1) <= fifo_full_139867185249696(0);
        
        fifo_inputs_139867185250200(3) <= outputs_139867185249752(2);
        outputs_full_139867185249752(2) <= fifo_full_139867185250200(3);
        
        fifo_inputs_139867185249304(2) <= outputs_139867185249752(3);
        outputs_full_139867185249752(3) <= fifo_full_139867185249304(2);
        
        fifo_inputs_139867185249864(1) <= outputs_139867185249808(0);
        outputs_full_139867185249808(0) <= fifo_full_139867185249864(1);
        
        fifo_inputs_139867185249752(0) <= outputs_139867185249808(1);
        outputs_full_139867185249808(1) <= fifo_full_139867185249752(0);
        
        fifo_inputs_139867185250256(3) <= outputs_139867185249808(2);
        outputs_full_139867185249808(2) <= fifo_full_139867185250256(3);
        
        fifo_inputs_139867185249360(2) <= outputs_139867185249808(3);
        outputs_full_139867185249808(3) <= fifo_full_139867185249360(2);
        
        fifo_inputs_139867185249920(1) <= outputs_139867185249864(0);
        outputs_full_139867185249864(0) <= fifo_full_139867185249920(1);
        
        fifo_inputs_139867185249808(0) <= outputs_139867185249864(1);
        outputs_full_139867185249864(1) <= fifo_full_139867185249808(0);
        
        fifo_inputs_139867185291336(3) <= outputs_139867185249864(2);
        outputs_full_139867185249864(2) <= fifo_full_139867185291336(3);
        
        fifo_inputs_139867185249416(2) <= outputs_139867185249864(3);
        outputs_full_139867185249864(3) <= fifo_full_139867185249416(2);
        
        fifo_inputs_139867185249976(1) <= outputs_139867185249920(0);
        outputs_full_139867185249920(0) <= fifo_full_139867185249976(1);
        
        fifo_inputs_139867185249864(0) <= outputs_139867185249920(1);
        outputs_full_139867185249920(1) <= fifo_full_139867185249864(0);
        
        fifo_inputs_139867185291392(3) <= outputs_139867185249920(2);
        outputs_full_139867185249920(2) <= fifo_full_139867185291392(3);
        
        fifo_inputs_139867185249472(2) <= outputs_139867185249920(3);
        outputs_full_139867185249920(3) <= fifo_full_139867185249472(2);
        
        fifo_inputs_139867185249920(0) <= outputs_139867185249976(1);
        outputs_full_139867185249976(1) <= fifo_full_139867185249920(0);
        
        fifo_inputs_139867185291448(3) <= outputs_139867185249976(2);
        outputs_full_139867185249976(2) <= fifo_full_139867185291448(3);
        
        fifo_inputs_139867185249528(2) <= outputs_139867185249976(3);
        outputs_full_139867185249976(3) <= fifo_full_139867185249528(2);
        
        fifo_inputs_139867185250088(1) <= outputs_139867185250032(0);
        outputs_full_139867185250032(0) <= fifo_full_139867185250088(1);
        
        fifo_inputs_139867185291504(3) <= outputs_139867185250032(2);
        outputs_full_139867185250032(2) <= fifo_full_139867185291504(3);
        
        fifo_inputs_139867185249584(2) <= outputs_139867185250032(3);
        outputs_full_139867185250032(3) <= fifo_full_139867185249584(2);
        
        fifo_inputs_139867185250144(1) <= outputs_139867185250088(0);
        outputs_full_139867185250088(0) <= fifo_full_139867185250144(1);
        
        fifo_inputs_139867185250032(0) <= outputs_139867185250088(1);
        outputs_full_139867185250088(1) <= fifo_full_139867185250032(0);
        
        fifo_inputs_139867185291560(3) <= outputs_139867185250088(2);
        outputs_full_139867185250088(2) <= fifo_full_139867185291560(3);
        
        fifo_inputs_139867185249640(2) <= outputs_139867185250088(3);
        outputs_full_139867185250088(3) <= fifo_full_139867185249640(2);
        
        fifo_inputs_139867185250200(1) <= outputs_139867185250144(0);
        outputs_full_139867185250144(0) <= fifo_full_139867185250200(1);
        
        fifo_inputs_139867185250088(0) <= outputs_139867185250144(1);
        outputs_full_139867185250144(1) <= fifo_full_139867185250088(0);
        
        fifo_inputs_139867185291616(3) <= outputs_139867185250144(2);
        outputs_full_139867185250144(2) <= fifo_full_139867185291616(3);
        
        fifo_inputs_139867185249696(2) <= outputs_139867185250144(3);
        outputs_full_139867185250144(3) <= fifo_full_139867185249696(2);
        
        fifo_inputs_139867185250256(1) <= outputs_139867185250200(0);
        outputs_full_139867185250200(0) <= fifo_full_139867185250256(1);
        
        fifo_inputs_139867185250144(0) <= outputs_139867185250200(1);
        outputs_full_139867185250200(1) <= fifo_full_139867185250144(0);
        
        fifo_inputs_139867185291672(3) <= outputs_139867185250200(2);
        outputs_full_139867185250200(2) <= fifo_full_139867185291672(3);
        
        fifo_inputs_139867185249752(2) <= outputs_139867185250200(3);
        outputs_full_139867185250200(3) <= fifo_full_139867185249752(2);
        
        fifo_inputs_139867185291336(1) <= outputs_139867185250256(0);
        outputs_full_139867185250256(0) <= fifo_full_139867185291336(1);
        
        fifo_inputs_139867185250200(0) <= outputs_139867185250256(1);
        outputs_full_139867185250256(1) <= fifo_full_139867185250200(0);
        
        fifo_inputs_139867185291728(3) <= outputs_139867185250256(2);
        outputs_full_139867185250256(2) <= fifo_full_139867185291728(3);
        
        fifo_inputs_139867185249808(2) <= outputs_139867185250256(3);
        outputs_full_139867185250256(3) <= fifo_full_139867185249808(2);
        
        fifo_inputs_139867185291392(1) <= outputs_139867185291336(0);
        outputs_full_139867185291336(0) <= fifo_full_139867185291392(1);
        
        fifo_inputs_139867185250256(0) <= outputs_139867185291336(1);
        outputs_full_139867185291336(1) <= fifo_full_139867185250256(0);
        
        fifo_inputs_139867185291784(3) <= outputs_139867185291336(2);
        outputs_full_139867185291336(2) <= fifo_full_139867185291784(3);
        
        fifo_inputs_139867185249864(2) <= outputs_139867185291336(3);
        outputs_full_139867185291336(3) <= fifo_full_139867185249864(2);
        
        fifo_inputs_139867185291448(1) <= outputs_139867185291392(0);
        outputs_full_139867185291392(0) <= fifo_full_139867185291448(1);
        
        fifo_inputs_139867185291336(0) <= outputs_139867185291392(1);
        outputs_full_139867185291392(1) <= fifo_full_139867185291336(0);
        
        fifo_inputs_139867185291840(3) <= outputs_139867185291392(2);
        outputs_full_139867185291392(2) <= fifo_full_139867185291840(3);
        
        fifo_inputs_139867185249920(2) <= outputs_139867185291392(3);
        outputs_full_139867185291392(3) <= fifo_full_139867185249920(2);
        
        fifo_inputs_139867185291392(0) <= outputs_139867185291448(1);
        outputs_full_139867185291448(1) <= fifo_full_139867185291392(0);
        
        fifo_inputs_139867185291896(3) <= outputs_139867185291448(2);
        outputs_full_139867185291448(2) <= fifo_full_139867185291896(3);
        
        fifo_inputs_139867185249976(2) <= outputs_139867185291448(3);
        outputs_full_139867185291448(3) <= fifo_full_139867185249976(2);
        
        fifo_inputs_139867185291560(1) <= outputs_139867185291504(0);
        outputs_full_139867185291504(0) <= fifo_full_139867185291560(1);
        
        fifo_inputs_139867185291952(3) <= outputs_139867185291504(2);
        outputs_full_139867185291504(2) <= fifo_full_139867185291952(3);
        
        fifo_inputs_139867185250032(2) <= outputs_139867185291504(3);
        outputs_full_139867185291504(3) <= fifo_full_139867185250032(2);
        
        fifo_inputs_139867185291616(1) <= outputs_139867185291560(0);
        outputs_full_139867185291560(0) <= fifo_full_139867185291616(1);
        
        fifo_inputs_139867185291504(0) <= outputs_139867185291560(1);
        outputs_full_139867185291560(1) <= fifo_full_139867185291504(0);
        
        fifo_inputs_139867185292008(3) <= outputs_139867185291560(2);
        outputs_full_139867185291560(2) <= fifo_full_139867185292008(3);
        
        fifo_inputs_139867185250088(2) <= outputs_139867185291560(3);
        outputs_full_139867185291560(3) <= fifo_full_139867185250088(2);
        
        fifo_inputs_139867185291672(1) <= outputs_139867185291616(0);
        outputs_full_139867185291616(0) <= fifo_full_139867185291672(1);
        
        fifo_inputs_139867185291560(0) <= outputs_139867185291616(1);
        outputs_full_139867185291616(1) <= fifo_full_139867185291560(0);
        
        fifo_inputs_139867185292064(3) <= outputs_139867185291616(2);
        outputs_full_139867185291616(2) <= fifo_full_139867185292064(3);
        
        fifo_inputs_139867185250144(2) <= outputs_139867185291616(3);
        outputs_full_139867185291616(3) <= fifo_full_139867185250144(2);
        
        fifo_inputs_139867185291728(1) <= outputs_139867185291672(0);
        outputs_full_139867185291672(0) <= fifo_full_139867185291728(1);
        
        fifo_inputs_139867185291616(0) <= outputs_139867185291672(1);
        outputs_full_139867185291672(1) <= fifo_full_139867185291616(0);
        
        fifo_inputs_139867185292120(3) <= outputs_139867185291672(2);
        outputs_full_139867185291672(2) <= fifo_full_139867185292120(3);
        
        fifo_inputs_139867185250200(2) <= outputs_139867185291672(3);
        outputs_full_139867185291672(3) <= fifo_full_139867185250200(2);
        
        fifo_inputs_139867185291784(1) <= outputs_139867185291728(0);
        outputs_full_139867185291728(0) <= fifo_full_139867185291784(1);
        
        fifo_inputs_139867185291672(0) <= outputs_139867185291728(1);
        outputs_full_139867185291728(1) <= fifo_full_139867185291672(0);
        
        fifo_inputs_139867185292176(3) <= outputs_139867185291728(2);
        outputs_full_139867185291728(2) <= fifo_full_139867185292176(3);
        
        fifo_inputs_139867185250256(2) <= outputs_139867185291728(3);
        outputs_full_139867185291728(3) <= fifo_full_139867185250256(2);
        
        fifo_inputs_139867185291840(1) <= outputs_139867185291784(0);
        outputs_full_139867185291784(0) <= fifo_full_139867185291840(1);
        
        fifo_inputs_139867185291728(0) <= outputs_139867185291784(1);
        outputs_full_139867185291784(1) <= fifo_full_139867185291728(0);
        
        fifo_inputs_139867185292232(3) <= outputs_139867185291784(2);
        outputs_full_139867185291784(2) <= fifo_full_139867185292232(3);
        
        fifo_inputs_139867185291336(2) <= outputs_139867185291784(3);
        outputs_full_139867185291784(3) <= fifo_full_139867185291336(2);
        
        fifo_inputs_139867185291896(1) <= outputs_139867185291840(0);
        outputs_full_139867185291840(0) <= fifo_full_139867185291896(1);
        
        fifo_inputs_139867185291784(0) <= outputs_139867185291840(1);
        outputs_full_139867185291840(1) <= fifo_full_139867185291784(0);
        
        fifo_inputs_139867185292288(3) <= outputs_139867185291840(2);
        outputs_full_139867185291840(2) <= fifo_full_139867185292288(3);
        
        fifo_inputs_139867185291392(2) <= outputs_139867185291840(3);
        outputs_full_139867185291840(3) <= fifo_full_139867185291392(2);
        
        fifo_inputs_139867185291840(0) <= outputs_139867185291896(1);
        outputs_full_139867185291896(1) <= fifo_full_139867185291840(0);
        
        fifo_inputs_139867185292344(3) <= outputs_139867185291896(2);
        outputs_full_139867185291896(2) <= fifo_full_139867185292344(3);
        
        fifo_inputs_139867185291448(2) <= outputs_139867185291896(3);
        outputs_full_139867185291896(3) <= fifo_full_139867185291448(2);
        
        fifo_inputs_139867185292008(1) <= outputs_139867185291952(0);
        outputs_full_139867185291952(0) <= fifo_full_139867185292008(1);
        
        fifo_inputs_139867185292400(3) <= outputs_139867185291952(2);
        outputs_full_139867185291952(2) <= fifo_full_139867185292400(3);
        
        fifo_inputs_139867185291504(2) <= outputs_139867185291952(3);
        outputs_full_139867185291952(3) <= fifo_full_139867185291504(2);
        
        fifo_inputs_139867185292064(1) <= outputs_139867185292008(0);
        outputs_full_139867185292008(0) <= fifo_full_139867185292064(1);
        
        fifo_inputs_139867185291952(0) <= outputs_139867185292008(1);
        outputs_full_139867185292008(1) <= fifo_full_139867185291952(0);
        
        fifo_inputs_139867185292456(3) <= outputs_139867185292008(2);
        outputs_full_139867185292008(2) <= fifo_full_139867185292456(3);
        
        fifo_inputs_139867185291560(2) <= outputs_139867185292008(3);
        outputs_full_139867185292008(3) <= fifo_full_139867185291560(2);
        
        fifo_inputs_139867185292120(1) <= outputs_139867185292064(0);
        outputs_full_139867185292064(0) <= fifo_full_139867185292120(1);
        
        fifo_inputs_139867185292008(0) <= outputs_139867185292064(1);
        outputs_full_139867185292064(1) <= fifo_full_139867185292008(0);
        
        fifo_inputs_139867185292512(3) <= outputs_139867185292064(2);
        outputs_full_139867185292064(2) <= fifo_full_139867185292512(3);
        
        fifo_inputs_139867185291616(2) <= outputs_139867185292064(3);
        outputs_full_139867185292064(3) <= fifo_full_139867185291616(2);
        
        fifo_inputs_139867185292176(1) <= outputs_139867185292120(0);
        outputs_full_139867185292120(0) <= fifo_full_139867185292176(1);
        
        fifo_inputs_139867185292064(0) <= outputs_139867185292120(1);
        outputs_full_139867185292120(1) <= fifo_full_139867185292064(0);
        
        fifo_inputs_139867185292568(3) <= outputs_139867185292120(2);
        outputs_full_139867185292120(2) <= fifo_full_139867185292568(3);
        
        fifo_inputs_139867185291672(2) <= outputs_139867185292120(3);
        outputs_full_139867185292120(3) <= fifo_full_139867185291672(2);
        
        fifo_inputs_139867185292232(1) <= outputs_139867185292176(0);
        outputs_full_139867185292176(0) <= fifo_full_139867185292232(1);
        
        fifo_inputs_139867185292120(0) <= outputs_139867185292176(1);
        outputs_full_139867185292176(1) <= fifo_full_139867185292120(0);
        
        fifo_inputs_139867185292624(3) <= outputs_139867185292176(2);
        outputs_full_139867185292176(2) <= fifo_full_139867185292624(3);
        
        fifo_inputs_139867185291728(2) <= outputs_139867185292176(3);
        outputs_full_139867185292176(3) <= fifo_full_139867185291728(2);
        
        fifo_inputs_139867185292288(1) <= outputs_139867185292232(0);
        outputs_full_139867185292232(0) <= fifo_full_139867185292288(1);
        
        fifo_inputs_139867185292176(0) <= outputs_139867185292232(1);
        outputs_full_139867185292232(1) <= fifo_full_139867185292176(0);
        
        fifo_inputs_139867185292680(3) <= outputs_139867185292232(2);
        outputs_full_139867185292232(2) <= fifo_full_139867185292680(3);
        
        fifo_inputs_139867185291784(2) <= outputs_139867185292232(3);
        outputs_full_139867185292232(3) <= fifo_full_139867185291784(2);
        
        fifo_inputs_139867185292344(1) <= outputs_139867185292288(0);
        outputs_full_139867185292288(0) <= fifo_full_139867185292344(1);
        
        fifo_inputs_139867185292232(0) <= outputs_139867185292288(1);
        outputs_full_139867185292288(1) <= fifo_full_139867185292232(0);
        
        fifo_inputs_139867185292736(3) <= outputs_139867185292288(2);
        outputs_full_139867185292288(2) <= fifo_full_139867185292736(3);
        
        fifo_inputs_139867185291840(2) <= outputs_139867185292288(3);
        outputs_full_139867185292288(3) <= fifo_full_139867185291840(2);
        
        fifo_inputs_139867185292288(0) <= outputs_139867185292344(1);
        outputs_full_139867185292344(1) <= fifo_full_139867185292288(0);
        
        fifo_inputs_139867185292792(3) <= outputs_139867185292344(2);
        outputs_full_139867185292344(2) <= fifo_full_139867185292792(3);
        
        fifo_inputs_139867185291896(2) <= outputs_139867185292344(3);
        outputs_full_139867185292344(3) <= fifo_full_139867185291896(2);
        
        fifo_inputs_139867185292456(1) <= outputs_139867185292400(0);
        outputs_full_139867185292400(0) <= fifo_full_139867185292456(1);
        
        fifo_inputs_139867185292848(3) <= outputs_139867185292400(2);
        outputs_full_139867185292400(2) <= fifo_full_139867185292848(3);
        
        fifo_inputs_139867185291952(2) <= outputs_139867185292400(3);
        outputs_full_139867185292400(3) <= fifo_full_139867185291952(2);
        
        fifo_inputs_139867185292512(1) <= outputs_139867185292456(0);
        outputs_full_139867185292456(0) <= fifo_full_139867185292512(1);
        
        fifo_inputs_139867185292400(0) <= outputs_139867185292456(1);
        outputs_full_139867185292456(1) <= fifo_full_139867185292400(0);
        
        fifo_inputs_139867185292904(3) <= outputs_139867185292456(2);
        outputs_full_139867185292456(2) <= fifo_full_139867185292904(3);
        
        fifo_inputs_139867185292008(2) <= outputs_139867185292456(3);
        outputs_full_139867185292456(3) <= fifo_full_139867185292008(2);
        
        fifo_inputs_139867185292568(1) <= outputs_139867185292512(0);
        outputs_full_139867185292512(0) <= fifo_full_139867185292568(1);
        
        fifo_inputs_139867185292456(0) <= outputs_139867185292512(1);
        outputs_full_139867185292512(1) <= fifo_full_139867185292456(0);
        
        fifo_inputs_139867185292960(3) <= outputs_139867185292512(2);
        outputs_full_139867185292512(2) <= fifo_full_139867185292960(3);
        
        fifo_inputs_139867185292064(2) <= outputs_139867185292512(3);
        outputs_full_139867185292512(3) <= fifo_full_139867185292064(2);
        
        fifo_inputs_139867185292624(1) <= outputs_139867185292568(0);
        outputs_full_139867185292568(0) <= fifo_full_139867185292624(1);
        
        fifo_inputs_139867185292512(0) <= outputs_139867185292568(1);
        outputs_full_139867185292568(1) <= fifo_full_139867185292512(0);
        
        fifo_inputs_139867185293016(3) <= outputs_139867185292568(2);
        outputs_full_139867185292568(2) <= fifo_full_139867185293016(3);
        
        fifo_inputs_139867185292120(2) <= outputs_139867185292568(3);
        outputs_full_139867185292568(3) <= fifo_full_139867185292120(2);
        
        fifo_inputs_139867185292680(1) <= outputs_139867185292624(0);
        outputs_full_139867185292624(0) <= fifo_full_139867185292680(1);
        
        fifo_inputs_139867185292568(0) <= outputs_139867185292624(1);
        outputs_full_139867185292624(1) <= fifo_full_139867185292568(0);
        
        fifo_inputs_139867185293072(3) <= outputs_139867185292624(2);
        outputs_full_139867185292624(2) <= fifo_full_139867185293072(3);
        
        fifo_inputs_139867185292176(2) <= outputs_139867185292624(3);
        outputs_full_139867185292624(3) <= fifo_full_139867185292176(2);
        
        fifo_inputs_139867185292736(1) <= outputs_139867185292680(0);
        outputs_full_139867185292680(0) <= fifo_full_139867185292736(1);
        
        fifo_inputs_139867185292624(0) <= outputs_139867185292680(1);
        outputs_full_139867185292680(1) <= fifo_full_139867185292624(0);
        
        fifo_inputs_139867185293128(3) <= outputs_139867185292680(2);
        outputs_full_139867185292680(2) <= fifo_full_139867185293128(3);
        
        fifo_inputs_139867185292232(2) <= outputs_139867185292680(3);
        outputs_full_139867185292680(3) <= fifo_full_139867185292232(2);
        
        fifo_inputs_139867185292792(1) <= outputs_139867185292736(0);
        outputs_full_139867185292736(0) <= fifo_full_139867185292792(1);
        
        fifo_inputs_139867185292680(0) <= outputs_139867185292736(1);
        outputs_full_139867185292736(1) <= fifo_full_139867185292680(0);
        
        fifo_inputs_139867185293184(3) <= outputs_139867185292736(2);
        outputs_full_139867185292736(2) <= fifo_full_139867185293184(3);
        
        fifo_inputs_139867185292288(2) <= outputs_139867185292736(3);
        outputs_full_139867185292736(3) <= fifo_full_139867185292288(2);
        
        fifo_inputs_139867185292736(0) <= outputs_139867185292792(1);
        outputs_full_139867185292792(1) <= fifo_full_139867185292736(0);
        
        fifo_inputs_139867185293240(3) <= outputs_139867185292792(2);
        outputs_full_139867185292792(2) <= fifo_full_139867185293240(3);
        
        fifo_inputs_139867185292344(2) <= outputs_139867185292792(3);
        outputs_full_139867185292792(3) <= fifo_full_139867185292344(2);
        
        fifo_inputs_139867185292904(1) <= outputs_139867185292848(0);
        outputs_full_139867185292848(0) <= fifo_full_139867185292904(1);
        
        fifo_inputs_139867185292400(2) <= outputs_139867185292848(3);
        outputs_full_139867185292848(3) <= fifo_full_139867185292400(2);
        
        fifo_inputs_139867185292960(1) <= outputs_139867185292904(0);
        outputs_full_139867185292904(0) <= fifo_full_139867185292960(1);
        
        fifo_inputs_139867185292848(0) <= outputs_139867185292904(1);
        outputs_full_139867185292904(1) <= fifo_full_139867185292848(0);
        
        fifo_inputs_139867185292456(2) <= outputs_139867185292904(3);
        outputs_full_139867185292904(3) <= fifo_full_139867185292456(2);
        
        fifo_inputs_139867185293016(1) <= outputs_139867185292960(0);
        outputs_full_139867185292960(0) <= fifo_full_139867185293016(1);
        
        fifo_inputs_139867185292904(0) <= outputs_139867185292960(1);
        outputs_full_139867185292960(1) <= fifo_full_139867185292904(0);
        
        fifo_inputs_139867185292512(2) <= outputs_139867185292960(3);
        outputs_full_139867185292960(3) <= fifo_full_139867185292512(2);
        
        fifo_inputs_139867185293072(1) <= outputs_139867185293016(0);
        outputs_full_139867185293016(0) <= fifo_full_139867185293072(1);
        
        fifo_inputs_139867185292960(0) <= outputs_139867185293016(1);
        outputs_full_139867185293016(1) <= fifo_full_139867185292960(0);
        
        fifo_inputs_139867185292568(2) <= outputs_139867185293016(3);
        outputs_full_139867185293016(3) <= fifo_full_139867185292568(2);
        
        fifo_inputs_139867185293128(1) <= outputs_139867185293072(0);
        outputs_full_139867185293072(0) <= fifo_full_139867185293128(1);
        
        fifo_inputs_139867185293016(0) <= outputs_139867185293072(1);
        outputs_full_139867185293072(1) <= fifo_full_139867185293016(0);
        
        fifo_inputs_139867185292624(2) <= outputs_139867185293072(3);
        outputs_full_139867185293072(3) <= fifo_full_139867185292624(2);
        
        fifo_inputs_139867185293184(1) <= outputs_139867185293128(0);
        outputs_full_139867185293128(0) <= fifo_full_139867185293184(1);
        
        fifo_inputs_139867185293072(0) <= outputs_139867185293128(1);
        outputs_full_139867185293128(1) <= fifo_full_139867185293072(0);
        
        fifo_inputs_139867185292680(2) <= outputs_139867185293128(3);
        outputs_full_139867185293128(3) <= fifo_full_139867185292680(2);
        
        fifo_inputs_139867185293240(1) <= outputs_139867185293184(0);
        outputs_full_139867185293184(0) <= fifo_full_139867185293240(1);
        
        fifo_inputs_139867185293128(0) <= outputs_139867185293184(1);
        outputs_full_139867185293184(1) <= fifo_full_139867185293128(0);
        
        fifo_inputs_139867185292736(2) <= outputs_139867185293184(3);
        outputs_full_139867185293184(3) <= fifo_full_139867185292736(2);
        
        fifo_inputs_139867185293184(0) <= outputs_139867185293240(1);
        outputs_full_139867185293240(1) <= fifo_full_139867185293184(0);
        
        fifo_inputs_139867185292792(2) <= outputs_139867185293240(3);
        outputs_full_139867185293240(3) <= fifo_full_139867185292792(2);
        

    
        core_inst_139867185248632: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185248632,
            fifo_full => fifo_full_139867185248632,
            outputs => outputs_139867185248632,
            outputs_full => outputs_full_139867185248632
        );
        
        core_inst_139867185248856: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185248856,
            fifo_full => fifo_full_139867185248856,
            outputs => outputs_139867185248856,
            outputs_full => outputs_full_139867185248856
        );
        
        core_inst_139867185248912: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185248912,
            fifo_full => fifo_full_139867185248912,
            outputs => outputs_139867185248912,
            outputs_full => outputs_full_139867185248912
        );
        
        core_inst_139867185248968: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185248968,
            fifo_full => fifo_full_139867185248968,
            outputs => outputs_139867185248968,
            outputs_full => outputs_full_139867185248968
        );
        
        core_inst_139867185248800: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185248800,
            fifo_full => fifo_full_139867185248800,
            outputs => outputs_139867185248800,
            outputs_full => outputs_full_139867185248800
        );
        
        core_inst_139867185249024: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185249024,
            fifo_full => fifo_full_139867185249024,
            outputs => outputs_139867185249024,
            outputs_full => outputs_full_139867185249024
        );
        
        core_inst_139867185249080: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185249080,
            fifo_full => fifo_full_139867185249080,
            outputs => outputs_139867185249080,
            outputs_full => outputs_full_139867185249080
        );
        
        core_inst_139867185249136: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185249136,
            fifo_full => fifo_full_139867185249136,
            outputs => outputs_139867185249136,
            outputs_full => outputs_full_139867185249136
        );
        
        core_inst_139867185249192: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185249192,
            fifo_full => fifo_full_139867185249192,
            outputs => outputs_139867185249192,
            outputs_full => outputs_full_139867185249192
        );
        
        core_inst_139867185248744: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185248744,
            fifo_full => fifo_full_139867185248744,
            outputs => outputs_139867185248744,
            outputs_full => outputs_full_139867185248744
        );
        
        core_inst_139867185249248: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185249248,
            fifo_full => fifo_full_139867185249248,
            outputs => outputs_139867185249248,
            outputs_full => outputs_full_139867185249248
        );
        
        core_inst_139867185249304: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185249304,
            fifo_full => fifo_full_139867185249304,
            outputs => outputs_139867185249304,
            outputs_full => outputs_full_139867185249304
        );
        
        core_inst_139867185249360: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185249360,
            fifo_full => fifo_full_139867185249360,
            outputs => outputs_139867185249360,
            outputs_full => outputs_full_139867185249360
        );
        
        core_inst_139867185249416: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185249416,
            fifo_full => fifo_full_139867185249416,
            outputs => outputs_139867185249416,
            outputs_full => outputs_full_139867185249416
        );
        
        core_inst_139867185249472: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185249472,
            fifo_full => fifo_full_139867185249472,
            outputs => outputs_139867185249472,
            outputs_full => outputs_full_139867185249472
        );
        
        core_inst_139867185249528: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185249528,
            fifo_full => fifo_full_139867185249528,
            outputs => outputs_139867185249528,
            outputs_full => outputs_full_139867185249528
        );
        
        core_inst_139867185249584: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185249584,
            fifo_full => fifo_full_139867185249584,
            outputs => outputs_139867185249584,
            outputs_full => outputs_full_139867185249584
        );
        
        core_inst_139867185249640: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185249640,
            fifo_full => fifo_full_139867185249640,
            outputs => outputs_139867185249640,
            outputs_full => outputs_full_139867185249640
        );
        
        core_inst_139867185249696: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185249696,
            fifo_full => fifo_full_139867185249696,
            outputs => outputs_139867185249696,
            outputs_full => outputs_full_139867185249696
        );
        
        core_inst_139867185249752: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185249752,
            fifo_full => fifo_full_139867185249752,
            outputs => outputs_139867185249752,
            outputs_full => outputs_full_139867185249752
        );
        
        core_inst_139867185249808: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185249808,
            fifo_full => fifo_full_139867185249808,
            outputs => outputs_139867185249808,
            outputs_full => outputs_full_139867185249808
        );
        
        core_inst_139867185249864: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185249864,
            fifo_full => fifo_full_139867185249864,
            outputs => outputs_139867185249864,
            outputs_full => outputs_full_139867185249864
        );
        
        core_inst_139867185249920: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185249920,
            fifo_full => fifo_full_139867185249920,
            outputs => outputs_139867185249920,
            outputs_full => outputs_full_139867185249920
        );
        
        core_inst_139867185249976: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185249976,
            fifo_full => fifo_full_139867185249976,
            outputs => outputs_139867185249976,
            outputs_full => outputs_full_139867185249976
        );
        
        core_inst_139867185250032: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185250032,
            fifo_full => fifo_full_139867185250032,
            outputs => outputs_139867185250032,
            outputs_full => outputs_full_139867185250032
        );
        
        core_inst_139867185250088: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185250088,
            fifo_full => fifo_full_139867185250088,
            outputs => outputs_139867185250088,
            outputs_full => outputs_full_139867185250088
        );
        
        core_inst_139867185250144: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185250144,
            fifo_full => fifo_full_139867185250144,
            outputs => outputs_139867185250144,
            outputs_full => outputs_full_139867185250144
        );
        
        core_inst_139867185250200: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185250200,
            fifo_full => fifo_full_139867185250200,
            outputs => outputs_139867185250200,
            outputs_full => outputs_full_139867185250200
        );
        
        core_inst_139867185250256: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185250256,
            fifo_full => fifo_full_139867185250256,
            outputs => outputs_139867185250256,
            outputs_full => outputs_full_139867185250256
        );
        
        core_inst_139867185291336: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185291336,
            fifo_full => fifo_full_139867185291336,
            outputs => outputs_139867185291336,
            outputs_full => outputs_full_139867185291336
        );
        
        core_inst_139867185291392: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185291392,
            fifo_full => fifo_full_139867185291392,
            outputs => outputs_139867185291392,
            outputs_full => outputs_full_139867185291392
        );
        
        core_inst_139867185291448: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185291448,
            fifo_full => fifo_full_139867185291448,
            outputs => outputs_139867185291448,
            outputs_full => outputs_full_139867185291448
        );
        
        core_inst_139867185291504: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185291504,
            fifo_full => fifo_full_139867185291504,
            outputs => outputs_139867185291504,
            outputs_full => outputs_full_139867185291504
        );
        
        core_inst_139867185291560: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185291560,
            fifo_full => fifo_full_139867185291560,
            outputs => outputs_139867185291560,
            outputs_full => outputs_full_139867185291560
        );
        
        core_inst_139867185291616: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185291616,
            fifo_full => fifo_full_139867185291616,
            outputs => outputs_139867185291616,
            outputs_full => outputs_full_139867185291616
        );
        
        core_inst_139867185291672: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185291672,
            fifo_full => fifo_full_139867185291672,
            outputs => outputs_139867185291672,
            outputs_full => outputs_full_139867185291672
        );
        
        core_inst_139867185291728: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185291728,
            fifo_full => fifo_full_139867185291728,
            outputs => outputs_139867185291728,
            outputs_full => outputs_full_139867185291728
        );
        
        core_inst_139867185291784: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185291784,
            fifo_full => fifo_full_139867185291784,
            outputs => outputs_139867185291784,
            outputs_full => outputs_full_139867185291784
        );
        
        core_inst_139867185291840: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185291840,
            fifo_full => fifo_full_139867185291840,
            outputs => outputs_139867185291840,
            outputs_full => outputs_full_139867185291840
        );
        
        core_inst_139867185291896: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185291896,
            fifo_full => fifo_full_139867185291896,
            outputs => outputs_139867185291896,
            outputs_full => outputs_full_139867185291896
        );
        
        core_inst_139867185291952: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185291952,
            fifo_full => fifo_full_139867185291952,
            outputs => outputs_139867185291952,
            outputs_full => outputs_full_139867185291952
        );
        
        core_inst_139867185292008: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185292008,
            fifo_full => fifo_full_139867185292008,
            outputs => outputs_139867185292008,
            outputs_full => outputs_full_139867185292008
        );
        
        core_inst_139867185292064: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185292064,
            fifo_full => fifo_full_139867185292064,
            outputs => outputs_139867185292064,
            outputs_full => outputs_full_139867185292064
        );
        
        core_inst_139867185292120: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185292120,
            fifo_full => fifo_full_139867185292120,
            outputs => outputs_139867185292120,
            outputs_full => outputs_full_139867185292120
        );
        
        core_inst_139867185292176: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185292176,
            fifo_full => fifo_full_139867185292176,
            outputs => outputs_139867185292176,
            outputs_full => outputs_full_139867185292176
        );
        
        core_inst_139867185292232: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185292232,
            fifo_full => fifo_full_139867185292232,
            outputs => outputs_139867185292232,
            outputs_full => outputs_full_139867185292232
        );
        
        core_inst_139867185292288: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185292288,
            fifo_full => fifo_full_139867185292288,
            outputs => outputs_139867185292288,
            outputs_full => outputs_full_139867185292288
        );
        
        core_inst_139867185292344: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185292344,
            fifo_full => fifo_full_139867185292344,
            outputs => outputs_139867185292344,
            outputs_full => outputs_full_139867185292344
        );
        
        core_inst_139867185292400: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185292400,
            fifo_full => fifo_full_139867185292400,
            outputs => outputs_139867185292400,
            outputs_full => outputs_full_139867185292400
        );
        
        core_inst_139867185292456: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185292456,
            fifo_full => fifo_full_139867185292456,
            outputs => outputs_139867185292456,
            outputs_full => outputs_full_139867185292456
        );
        
        core_inst_139867185292512: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185292512,
            fifo_full => fifo_full_139867185292512,
            outputs => outputs_139867185292512,
            outputs_full => outputs_full_139867185292512
        );
        
        core_inst_139867185292568: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185292568,
            fifo_full => fifo_full_139867185292568,
            outputs => outputs_139867185292568,
            outputs_full => outputs_full_139867185292568
        );
        
        core_inst_139867185292624: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185292624,
            fifo_full => fifo_full_139867185292624,
            outputs => outputs_139867185292624,
            outputs_full => outputs_full_139867185292624
        );
        
        core_inst_139867185292680: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185292680,
            fifo_full => fifo_full_139867185292680,
            outputs => outputs_139867185292680,
            outputs_full => outputs_full_139867185292680
        );
        
        core_inst_139867185292736: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185292736,
            fifo_full => fifo_full_139867185292736,
            outputs => outputs_139867185292736,
            outputs_full => outputs_full_139867185292736
        );
        
        core_inst_139867185292792: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185292792,
            fifo_full => fifo_full_139867185292792,
            outputs => outputs_139867185292792,
            outputs_full => outputs_full_139867185292792
        );
        
        core_inst_139867185292848: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185292848,
            fifo_full => fifo_full_139867185292848,
            outputs => outputs_139867185292848,
            outputs_full => outputs_full_139867185292848
        );
        
        core_inst_139867185292904: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185292904,
            fifo_full => fifo_full_139867185292904,
            outputs => outputs_139867185292904,
            outputs_full => outputs_full_139867185292904
        );
        
        core_inst_139867185292960: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185292960,
            fifo_full => fifo_full_139867185292960,
            outputs => outputs_139867185292960,
            outputs_full => outputs_full_139867185292960
        );
        
        core_inst_139867185293016: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185293016,
            fifo_full => fifo_full_139867185293016,
            outputs => outputs_139867185293016,
            outputs_full => outputs_full_139867185293016
        );
        
        core_inst_139867185293072: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185293072,
            fifo_full => fifo_full_139867185293072,
            outputs => outputs_139867185293072,
            outputs_full => outputs_full_139867185293072
        );
        
        core_inst_139867185293128: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185293128,
            fifo_full => fifo_full_139867185293128,
            outputs => outputs_139867185293128,
            outputs_full => outputs_full_139867185293128
        );
        
        core_inst_139867185293184: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185293184,
            fifo_full => fifo_full_139867185293184,
            outputs => outputs_139867185293184,
            outputs_full => outputs_full_139867185293184
        );
        
        core_inst_139867185293240: entity Core
        port map (
            clk => clk,
            clk_en => clk_en,
            reset => reset,
            addr => addr,
            data => data,
            we => we,
            fifo_inputs => fifo_inputs_139867185293240,
            fifo_full => fifo_full_139867185293240,
            outputs => outputs_139867185293240,
            outputs_full => outputs_full_139867185293240
        );
        

end behav;

